module matrix_adc_pipe (
    input         clk,
	input         rst, // High_active

    // INPUT DATA
    input  [159:0] in_dat,
	
	// COE DATA
	input  [159:0] coe_dat00, coe_dat01, coe_dat02, coe_dat03, coe_dat04, coe_dat05, coe_dat06,
                   coe_dat07, coe_dat08, coe_dat09, coe_dat10, coe_dat11, coe_dat12,
                   coe_dat13, coe_dat14, coe_dat15, coe_dat16, coe_dat17, coe_dat18,
                   coe_dat19, coe_dat20, coe_dat21, coe_dat22, coe_dat23, coe_dat24,
                   coe_dat25, coe_dat26, coe_dat27, coe_dat28, coe_dat29, coe_dat30, coe_dat31,
	input          loop_flg,
    input    [3:0] STATE,
	input    [5:0] cyc32_cnt,
    input    [4:0] row1_cnt,
	output         out_en,
	output  [19:0] out_dat
);

    parameter DLY=0.1;
    parameter ST_IDLE=4'd0;
	parameter ST_LOAD=4'd1;
	parameter ST_LOAD2=4'd2;
	parameter ST_EXEC=4'd3;
	parameter ST_JUDGE=4'd4;
	
//**********************************************************
//**********************************************************
	// PIPELINE
    reg [41:0]  pipeline_cnt ;
	reg [41:0]  loop_flg_hld ;
    reg [159:0] in_dat_dd1,  in_dat_dd2,  in_dat_dd3,  in_dat_dd4,
                in_dat_dd5,  in_dat_dd6,  in_dat_dd7,  in_dat_dd8,
                in_dat_dd9,  in_dat_dd10, in_dat_dd11, in_dat_dd12,
                in_dat_dd13, in_dat_dd14, in_dat_dd15, in_dat_dd16,
                in_dat_dd17, in_dat_dd18, in_dat_dd19, in_dat_dd20,
                in_dat_dd21, in_dat_dd22, in_dat_dd23, in_dat_dd24,
                in_dat_dd25, in_dat_dd26, in_dat_dd27, in_dat_dd28,
                in_dat_dd29, in_dat_dd30, in_dat_dd31, in_dat_dd32;
    reg [159:0] coe_dat00_dd, coe_dat01_dd, coe_dat02_dd, coe_dat03_dd,
                coe_dat04_dd, coe_dat05_dd, coe_dat06_dd, coe_dat07_dd,
                coe_dat08_dd, coe_dat09_dd, coe_dat10_dd, coe_dat11_dd,
                coe_dat12_dd, coe_dat13_dd, coe_dat14_dd, coe_dat15_dd,
                coe_dat16_dd, coe_dat17_dd, coe_dat18_dd, coe_dat19_dd,
                coe_dat20_dd, coe_dat21_dd, coe_dat22_dd, coe_dat23_dd,
                coe_dat24_dd, coe_dat25_dd, coe_dat26_dd, coe_dat27_dd,
                coe_dat28_dd, coe_dat29_dd, coe_dat30_dd, coe_dat31_dd;
 
    reg [5:0] cyc32_cnt_dd0,  cyc32_cnt_dd1,  cyc32_cnt_dd2,  cyc32_cnt_dd3,  cyc32_cnt_dd4,
              cyc32_cnt_dd5,  cyc32_cnt_dd6,  cyc32_cnt_dd7,  cyc32_cnt_dd8,  cyc32_cnt_dd9,
              cyc32_cnt_dd10, cyc32_cnt_dd11, cyc32_cnt_dd12, cyc32_cnt_dd13, cyc32_cnt_dd14,
              cyc32_cnt_dd15, cyc32_cnt_dd16, cyc32_cnt_dd17, cyc32_cnt_dd18, cyc32_cnt_dd19,
              cyc32_cnt_dd20, cyc32_cnt_dd21, cyc32_cnt_dd22, cyc32_cnt_dd23, cyc32_cnt_dd24,
              cyc32_cnt_dd25, cyc32_cnt_dd26, cyc32_cnt_dd27, cyc32_cnt_dd28, cyc32_cnt_dd29,
              cyc32_cnt_dd30, cyc32_cnt_dd31, cyc32_cnt_dd32, cyc32_cnt_dd33, cyc32_cnt_dd34,
              cyc32_cnt_dd35, cyc32_cnt_dd36, cyc32_cnt_dd37, cyc32_cnt_dd38, cyc32_cnt_dd39,
              cyc32_cnt_dd40, cyc32_cnt_dd41, cyc32_cnt_dd42;
	                       
                           
    always @ (posedge clk) begin
		if(rst) begin
		    cyc32_cnt_dd0[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd1[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd2[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd3[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd4[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd5[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd6[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd7[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd8[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd9[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd10[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd11[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd12[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd13[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd14[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd15[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd16[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd17[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd18[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd19[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd20[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd21[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd22[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd23[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd24[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd25[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd26[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd27[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd28[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd29[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd30[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd31[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd32[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd33[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd34[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd35[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd36[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd37[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd38[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd39[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd40[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd41[5:0] <= #DLY 6'd0 ;
		    cyc32_cnt_dd42[5:0] <= #DLY 6'd0 ;
		end else begin
		    cyc32_cnt_dd0[5:0]  <= #DLY cyc32_cnt[5:0] ;
		    cyc32_cnt_dd1[5:0]  <= #DLY cyc32_cnt_dd0[5:0] ;
		    cyc32_cnt_dd2[5:0]  <= #DLY cyc32_cnt_dd1[5:0] ;
		    cyc32_cnt_dd3[5:0]  <= #DLY cyc32_cnt_dd2[5:0] ;
		    cyc32_cnt_dd4[5:0]  <= #DLY cyc32_cnt_dd3[5:0] ;
		    cyc32_cnt_dd5[5:0]  <= #DLY cyc32_cnt_dd4[5:0] ;
		    cyc32_cnt_dd6[5:0]  <= #DLY cyc32_cnt_dd5[5:0] ;
		    cyc32_cnt_dd7[5:0]  <= #DLY cyc32_cnt_dd6[5:0] ;
		    cyc32_cnt_dd8[5:0]  <= #DLY cyc32_cnt_dd7[5:0] ;
		    cyc32_cnt_dd9[5:0]  <= #DLY cyc32_cnt_dd8[5:0] ;
		    cyc32_cnt_dd10[5:0] <= #DLY cyc32_cnt_dd9[5:0] ;
		    cyc32_cnt_dd11[5:0] <= #DLY cyc32_cnt_dd10[5:0] ;
		    cyc32_cnt_dd12[5:0] <= #DLY cyc32_cnt_dd11[5:0] ;
		    cyc32_cnt_dd13[5:0] <= #DLY cyc32_cnt_dd12[5:0] ;
		    cyc32_cnt_dd14[5:0] <= #DLY cyc32_cnt_dd13[5:0] ;
		    cyc32_cnt_dd15[5:0] <= #DLY cyc32_cnt_dd14[5:0] ;
		    cyc32_cnt_dd16[5:0] <= #DLY cyc32_cnt_dd15[5:0] ;
		    cyc32_cnt_dd17[5:0] <= #DLY cyc32_cnt_dd16[5:0] ;
		    cyc32_cnt_dd18[5:0] <= #DLY cyc32_cnt_dd17[5:0] ;
		    cyc32_cnt_dd19[5:0] <= #DLY cyc32_cnt_dd18[5:0] ;
		    cyc32_cnt_dd20[5:0] <= #DLY cyc32_cnt_dd19[5:0] ;
		    cyc32_cnt_dd21[5:0] <= #DLY cyc32_cnt_dd20[5:0] ;
		    cyc32_cnt_dd22[5:0] <= #DLY cyc32_cnt_dd21[5:0] ;
		    cyc32_cnt_dd23[5:0] <= #DLY cyc32_cnt_dd22[5:0] ;
		    cyc32_cnt_dd24[5:0] <= #DLY cyc32_cnt_dd23[5:0] ;
		    cyc32_cnt_dd25[5:0] <= #DLY cyc32_cnt_dd24[5:0] ;
		    cyc32_cnt_dd26[5:0] <= #DLY cyc32_cnt_dd25[5:0] ;
		    cyc32_cnt_dd27[5:0] <= #DLY cyc32_cnt_dd26[5:0] ;
		    cyc32_cnt_dd28[5:0] <= #DLY cyc32_cnt_dd27[5:0] ;
		    cyc32_cnt_dd29[5:0] <= #DLY cyc32_cnt_dd28[5:0] ;
		    cyc32_cnt_dd30[5:0] <= #DLY cyc32_cnt_dd29[5:0] ;
		    cyc32_cnt_dd31[5:0] <= #DLY cyc32_cnt_dd30[5:0] ;
		    cyc32_cnt_dd32[5:0] <= #DLY cyc32_cnt_dd31[5:0] ;
		    cyc32_cnt_dd33[5:0] <= #DLY cyc32_cnt_dd32[5:0] ;
		    cyc32_cnt_dd34[5:0] <= #DLY cyc32_cnt_dd33[5:0] ;
		    cyc32_cnt_dd35[5:0] <= #DLY cyc32_cnt_dd34[5:0] ;
		    cyc32_cnt_dd36[5:0] <= #DLY cyc32_cnt_dd35[5:0] ;
		    cyc32_cnt_dd37[5:0] <= #DLY cyc32_cnt_dd36[5:0] ;
		    cyc32_cnt_dd38[5:0] <= #DLY cyc32_cnt_dd37[5:0] ;
		    cyc32_cnt_dd39[5:0] <= #DLY cyc32_cnt_dd38[5:0] ;
		    cyc32_cnt_dd40[5:0] <= #DLY cyc32_cnt_dd39[5:0] ;
		    cyc32_cnt_dd41[5:0] <= #DLY cyc32_cnt_dd40[5:0] ;
		    cyc32_cnt_dd42[5:0] <= #DLY cyc32_cnt_dd41[5:0] ;
		end
	end


    always @ (posedge clk) begin
		if(rst) begin
            pipeline_cnt[41:0] <= #DLY 42'd0 ;
            loop_flg_hld[41:0] <= #DLY 42'd0 ;
		end else begin
            pipeline_cnt[41:0] <= #DLY {pipeline_cnt[40:0], (STATE[3:0]==ST_LOAD)} ;
            loop_flg_hld[41:0] <= #DLY {loop_flg_hld[40:0], (loop_flg & (STATE[3:0]==ST_LOAD))} ;
		end
	end

    always @ (posedge clk) begin
		if(rst) begin
			in_dat_dd1[159:0]  <= #DLY 160'd0 ;
			in_dat_dd2[159:0]  <= #DLY 160'd0 ;
			in_dat_dd3[159:0]  <= #DLY 160'd0 ;
			in_dat_dd4[159:0]  <= #DLY 160'd0 ;
			in_dat_dd5[159:0]  <= #DLY 160'd0 ;
			in_dat_dd6[159:0]  <= #DLY 160'd0 ;
			in_dat_dd7[159:0]  <= #DLY 160'd0 ;
			in_dat_dd8[159:0]  <= #DLY 160'd0 ;
			in_dat_dd9[159:0]  <= #DLY 160'd0 ;
			in_dat_dd10[159:0] <= #DLY 160'd0 ;
			in_dat_dd11[159:0] <= #DLY 160'd0 ;
			in_dat_dd12[159:0] <= #DLY 160'd0 ;
			in_dat_dd13[159:0] <= #DLY 160'd0 ;
			in_dat_dd14[159:0] <= #DLY 160'd0 ;
			in_dat_dd15[159:0] <= #DLY 160'd0 ;
			in_dat_dd16[159:0] <= #DLY 160'd0 ;
			in_dat_dd17[159:0] <= #DLY 160'd0 ;
			in_dat_dd18[159:0] <= #DLY 160'd0 ;
			in_dat_dd19[159:0] <= #DLY 160'd0 ;
			in_dat_dd20[159:0] <= #DLY 160'd0 ;
			in_dat_dd21[159:0] <= #DLY 160'd0 ;
			in_dat_dd22[159:0] <= #DLY 160'd0 ;
			in_dat_dd23[159:0] <= #DLY 160'd0 ;
			in_dat_dd24[159:0] <= #DLY 160'd0 ;
			in_dat_dd25[159:0] <= #DLY 160'd0 ;
			in_dat_dd26[159:0] <= #DLY 160'd0 ;
			in_dat_dd27[159:0] <= #DLY 160'd0 ;
			in_dat_dd28[159:0] <= #DLY 160'd0 ;
			in_dat_dd29[159:0] <= #DLY 160'd0 ;
			in_dat_dd30[159:0] <= #DLY 160'd0 ;
			in_dat_dd31[159:0] <= #DLY 160'd0 ;
			in_dat_dd32[159:0] <= #DLY 160'd0 ;
			
			coe_dat00_dd[159:0] <= #DLY 160'd0 ;
			coe_dat01_dd[159:0] <= #DLY 160'd0 ;
			coe_dat02_dd[159:0] <= #DLY 160'd0 ;
			coe_dat03_dd[159:0] <= #DLY 160'd0 ;
			coe_dat04_dd[159:0] <= #DLY 160'd0 ;
			coe_dat05_dd[159:0] <= #DLY 160'd0 ;
			coe_dat06_dd[159:0] <= #DLY 160'd0 ;
			coe_dat07_dd[159:0] <= #DLY 160'd0 ;
			coe_dat08_dd[159:0] <= #DLY 160'd0 ;
			coe_dat09_dd[159:0] <= #DLY 160'd0 ;
			coe_dat10_dd[159:0] <= #DLY 160'd0 ;
			coe_dat11_dd[159:0] <= #DLY 160'd0 ;
			coe_dat12_dd[159:0] <= #DLY 160'd0 ;
			coe_dat13_dd[159:0] <= #DLY 160'd0 ;
			coe_dat14_dd[159:0] <= #DLY 160'd0 ;
			coe_dat15_dd[159:0] <= #DLY 160'd0 ;
			coe_dat16_dd[159:0] <= #DLY 160'd0 ;
			coe_dat17_dd[159:0] <= #DLY 160'd0 ;
			coe_dat18_dd[159:0] <= #DLY 160'd0 ;
			coe_dat19_dd[159:0] <= #DLY 160'd0 ;
			coe_dat20_dd[159:0] <= #DLY 160'd0 ;
			coe_dat21_dd[159:0] <= #DLY 160'd0 ;
			coe_dat22_dd[159:0] <= #DLY 160'd0 ;
			coe_dat23_dd[159:0] <= #DLY 160'd0 ;
			coe_dat24_dd[159:0] <= #DLY 160'd0 ;
			coe_dat25_dd[159:0] <= #DLY 160'd0 ;
			coe_dat26_dd[159:0] <= #DLY 160'd0 ;
			coe_dat27_dd[159:0] <= #DLY 160'd0 ;
			coe_dat28_dd[159:0] <= #DLY 160'd0 ;
			coe_dat29_dd[159:0] <= #DLY 160'd0 ;
			coe_dat30_dd[159:0] <= #DLY 160'd0 ;
			coe_dat31_dd[159:0] <= #DLY 160'd0 ;			
		end else begin
            coe_dat00_dd[159:0] <= #DLY coe_dat00[159:0] ;
            coe_dat01_dd[159:0] <= #DLY coe_dat01[159:0] ;
            coe_dat02_dd[159:0] <= #DLY coe_dat02[159:0] ;
            coe_dat03_dd[159:0] <= #DLY coe_dat03[159:0] ;
            coe_dat04_dd[159:0] <= #DLY coe_dat04[159:0] ;
            coe_dat05_dd[159:0] <= #DLY coe_dat05[159:0] ;
            coe_dat06_dd[159:0] <= #DLY coe_dat06[159:0] ;
            coe_dat07_dd[159:0] <= #DLY coe_dat07[159:0] ;
            coe_dat08_dd[159:0] <= #DLY coe_dat08[159:0] ;
            coe_dat09_dd[159:0] <= #DLY coe_dat09[159:0] ;
            coe_dat10_dd[159:0] <= #DLY coe_dat10[159:0] ;
            coe_dat11_dd[159:0] <= #DLY coe_dat11[159:0] ;
            coe_dat12_dd[159:0] <= #DLY coe_dat12[159:0] ;
            coe_dat13_dd[159:0] <= #DLY coe_dat13[159:0] ;
            coe_dat14_dd[159:0] <= #DLY coe_dat14[159:0] ;
            coe_dat15_dd[159:0] <= #DLY coe_dat15[159:0] ;
            coe_dat16_dd[159:0] <= #DLY coe_dat16[159:0] ;
            coe_dat17_dd[159:0] <= #DLY coe_dat17[159:0] ;
            coe_dat18_dd[159:0] <= #DLY coe_dat18[159:0] ;
            coe_dat19_dd[159:0] <= #DLY coe_dat19[159:0] ;
            coe_dat20_dd[159:0] <= #DLY coe_dat20[159:0] ;
            coe_dat21_dd[159:0] <= #DLY coe_dat21[159:0] ;
            coe_dat22_dd[159:0] <= #DLY coe_dat22[159:0] ;
            coe_dat23_dd[159:0] <= #DLY coe_dat23[159:0] ;
            coe_dat24_dd[159:0] <= #DLY coe_dat24[159:0] ;
            coe_dat25_dd[159:0] <= #DLY coe_dat25[159:0] ;
            coe_dat26_dd[159:0] <= #DLY coe_dat26[159:0] ;
            coe_dat27_dd[159:0] <= #DLY coe_dat27[159:0] ;
            coe_dat28_dd[159:0] <= #DLY coe_dat28[159:0] ;
            coe_dat29_dd[159:0] <= #DLY coe_dat29[159:0] ;
            coe_dat30_dd[159:0] <= #DLY coe_dat30[159:0] ;
            coe_dat31_dd[159:0] <= #DLY coe_dat31[159:0] ;
			
			if(pipeline_cnt[0]) begin
				in_dat_dd1[159:0]  <= #DLY in_dat[159:0]      ;
				in_dat_dd2[159:0]  <= #DLY in_dat_dd1[159:0]  ;
				in_dat_dd3[159:0]  <= #DLY in_dat_dd2[159:0]  ;
				in_dat_dd4[159:0]  <= #DLY in_dat_dd3[159:0]  ;
				in_dat_dd5[159:0]  <= #DLY in_dat_dd4[159:0]  ;
				in_dat_dd6[159:0]  <= #DLY in_dat_dd5[159:0]  ;
				in_dat_dd7[159:0]  <= #DLY in_dat_dd6[159:0]  ;
				in_dat_dd8[159:0]  <= #DLY in_dat_dd7[159:0]  ;
				in_dat_dd9[159:0]  <= #DLY in_dat_dd8[159:0]  ;
				in_dat_dd10[159:0] <= #DLY in_dat_dd9[159:0]  ;
				in_dat_dd11[159:0] <= #DLY in_dat_dd10[159:0] ;
				in_dat_dd12[159:0] <= #DLY in_dat_dd11[159:0] ;
				in_dat_dd13[159:0] <= #DLY in_dat_dd12[159:0] ;
				in_dat_dd14[159:0] <= #DLY in_dat_dd13[159:0] ;
				in_dat_dd15[159:0] <= #DLY in_dat_dd14[159:0] ;
				in_dat_dd16[159:0] <= #DLY in_dat_dd15[159:0] ;
				in_dat_dd17[159:0] <= #DLY in_dat_dd16[159:0] ;
				in_dat_dd18[159:0] <= #DLY in_dat_dd17[159:0] ;
				in_dat_dd19[159:0] <= #DLY in_dat_dd18[159:0] ;
				in_dat_dd20[159:0] <= #DLY in_dat_dd19[159:0] ;
				in_dat_dd21[159:0] <= #DLY in_dat_dd20[159:0] ;
				in_dat_dd22[159:0] <= #DLY in_dat_dd21[159:0] ;
				in_dat_dd23[159:0] <= #DLY in_dat_dd22[159:0] ;
				in_dat_dd24[159:0] <= #DLY in_dat_dd23[159:0] ;
				in_dat_dd25[159:0] <= #DLY in_dat_dd24[159:0] ;
				in_dat_dd26[159:0] <= #DLY in_dat_dd25[159:0] ;
				in_dat_dd27[159:0] <= #DLY in_dat_dd26[159:0] ;
				in_dat_dd28[159:0] <= #DLY in_dat_dd27[159:0] ;
				in_dat_dd29[159:0] <= #DLY in_dat_dd28[159:0] ;
				in_dat_dd30[159:0] <= #DLY in_dat_dd29[159:0] ;
				in_dat_dd31[159:0] <= #DLY in_dat_dd30[159:0] ;
				in_dat_dd32[159:0] <= #DLY in_dat_dd31[159:0] ;
			end
		end
	end

///////////////////////////////////////////
// pipeline_cnt[] active
///////////////////////////////////////////


    wire [5119:0] in_dat_wire  = {in_dat_dd32[159:0], in_dat_dd31[159:0], in_dat_dd30[159:0], in_dat_dd29[159:0],
	                              in_dat_dd28[159:0], in_dat_dd27[159:0], in_dat_dd26[159:0], in_dat_dd25[159:0], 
	                              in_dat_dd24[159:0], in_dat_dd23[159:0], in_dat_dd22[159:0], in_dat_dd21[159:0], 
	                              in_dat_dd20[159:0], in_dat_dd19[159:0], in_dat_dd18[159:0], in_dat_dd17[159:0], 
	                              in_dat_dd16[159:0], in_dat_dd15[159:0], in_dat_dd14[159:0], in_dat_dd13[159:0], 
	                              in_dat_dd12[159:0], in_dat_dd11[159:0], in_dat_dd10[159:0], in_dat_dd9[159:0], 
	                              in_dat_dd8[159:0],  in_dat_dd7[159:0],  in_dat_dd6[159:0],  in_dat_dd5[159:0], 
	                              in_dat_dd4[159:0],  in_dat_dd3[159:0],  in_dat_dd2[159:0],  in_dat_dd1[159:0]};

    wire [5119:0] coe_dat_wire  = {coe_dat00[159:0], coe_dat01[159:0], coe_dat02[159:0], coe_dat03[159:0],
	                               coe_dat04[159:0], coe_dat05[159:0], coe_dat06[159:0], coe_dat07[159:0],
								   coe_dat08[159:0], coe_dat09[159:0], coe_dat10[159:0], coe_dat11[159:0],
								   coe_dat12[159:0], coe_dat13[159:0], coe_dat14[159:0], coe_dat15[159:0],
								   coe_dat16[159:0], coe_dat17[159:0], coe_dat18[159:0], coe_dat19[159:0],
								   coe_dat20[159:0], coe_dat21[159:0], coe_dat22[159:0], coe_dat23[159:0],
								   coe_dat24[159:0], coe_dat25[159:0], coe_dat26[159:0], coe_dat27[159:0],
								   coe_dat28[159:0], coe_dat29[159:0], coe_dat30[159:0], coe_dat31[159:0]};

    wire [9:0] in_dat_wire01  = in_dat_wire[5119:5110] ;
    wire [9:0] in_dat_wire02  = in_dat_wire[5109:5100] ;
    wire [9:0] in_dat_wire03  = in_dat_wire[5099:5090] ;
    wire [9:0] in_dat_wire04  = in_dat_wire[5089:5080] ;
    wire [9:0] in_dat_wire05  = in_dat_wire[5079:5070] ;
    wire [9:0] in_dat_wire06  = in_dat_wire[5069:5060] ;
    wire [9:0] in_dat_wire07  = in_dat_wire[5059:5050] ;
    wire [9:0] in_dat_wire08  = in_dat_wire[5049:5040] ;
    wire [9:0] in_dat_wire09  = in_dat_wire[5039:5030] ;
    wire [9:0] in_dat_wire10  = in_dat_wire[5029:5020] ;
    wire [9:0] in_dat_wire11  = in_dat_wire[5019:5010] ;
    wire [9:0] in_dat_wire12  = in_dat_wire[5009:5000] ;
    wire [9:0] in_dat_wire13  = in_dat_wire[4999:4990] ;
    wire [9:0] in_dat_wire14  = in_dat_wire[4989:4980] ;
    wire [9:0] in_dat_wire15  = in_dat_wire[4979:4970] ;
    wire [9:0] in_dat_wire16  = in_dat_wire[4969:4960] ;
    wire [9:0] in_dat_wire17  = in_dat_wire[4959:4950] ;
    wire [9:0] in_dat_wire18  = in_dat_wire[4949:4940] ;
    wire [9:0] in_dat_wire19  = in_dat_wire[4939:4930] ;
    wire [9:0] in_dat_wire20  = in_dat_wire[4929:4920] ;
    wire [9:0] in_dat_wire21  = in_dat_wire[4919:4910] ;
    wire [9:0] in_dat_wire22  = in_dat_wire[4909:4900] ;
    wire [9:0] in_dat_wire23  = in_dat_wire[4899:4890] ;
    wire [9:0] in_dat_wire24  = in_dat_wire[4889:4880] ;
    wire [9:0] in_dat_wire25  = in_dat_wire[4879:4870] ;
    wire [9:0] in_dat_wire26  = in_dat_wire[4869:4860] ;
    wire [9:0] in_dat_wire27  = in_dat_wire[4859:4850] ;
    wire [9:0] in_dat_wire28  = in_dat_wire[4849:4840] ;
    wire [9:0] in_dat_wire29  = in_dat_wire[4839:4830] ;
    wire [9:0] in_dat_wire30  = in_dat_wire[4829:4820] ;
    wire [9:0] in_dat_wire31  = in_dat_wire[4819:4810] ;
    wire [9:0] in_dat_wire32  = in_dat_wire[4809:4800] ;
    wire [9:0] in_dat_wire33  = in_dat_wire[4799:4790] ;
    wire [9:0] in_dat_wire34  = in_dat_wire[4789:4780] ;
    wire [9:0] in_dat_wire35  = in_dat_wire[4779:4770] ;
    wire [9:0] in_dat_wire36  = in_dat_wire[4769:4760] ;
    wire [9:0] in_dat_wire37  = in_dat_wire[4759:4750] ;
    wire [9:0] in_dat_wire38  = in_dat_wire[4749:4740] ;
    wire [9:0] in_dat_wire39  = in_dat_wire[4739:4730] ;
    wire [9:0] in_dat_wire40  = in_dat_wire[4729:4720] ;
    wire [9:0] in_dat_wire41  = in_dat_wire[4719:4710] ;
    wire [9:0] in_dat_wire42  = in_dat_wire[4709:4700] ;
    wire [9:0] in_dat_wire43  = in_dat_wire[4699:4690] ;
    wire [9:0] in_dat_wire44  = in_dat_wire[4689:4680] ;
    wire [9:0] in_dat_wire45  = in_dat_wire[4679:4670] ;
    wire [9:0] in_dat_wire46  = in_dat_wire[4669:4660] ;
    wire [9:0] in_dat_wire47  = in_dat_wire[4659:4650] ;
    wire [9:0] in_dat_wire48  = in_dat_wire[4649:4640] ;
    wire [9:0] in_dat_wire49  = in_dat_wire[4639:4630] ;
    wire [9:0] in_dat_wire50  = in_dat_wire[4629:4620] ;
    wire [9:0] in_dat_wire51  = in_dat_wire[4619:4610] ;
    wire [9:0] in_dat_wire52  = in_dat_wire[4609:4600] ;
    wire [9:0] in_dat_wire53  = in_dat_wire[4599:4590] ;
    wire [9:0] in_dat_wire54  = in_dat_wire[4589:4580] ;
    wire [9:0] in_dat_wire55  = in_dat_wire[4579:4570] ;
    wire [9:0] in_dat_wire56  = in_dat_wire[4569:4560] ;
    wire [9:0] in_dat_wire57  = in_dat_wire[4559:4550] ;
    wire [9:0] in_dat_wire58  = in_dat_wire[4549:4540] ;
    wire [9:0] in_dat_wire59  = in_dat_wire[4539:4530] ;
    wire [9:0] in_dat_wire60  = in_dat_wire[4529:4520] ;
    wire [9:0] in_dat_wire61  = in_dat_wire[4519:4510] ;
    wire [9:0] in_dat_wire62  = in_dat_wire[4509:4500] ;
    wire [9:0] in_dat_wire63  = in_dat_wire[4499:4490] ;
    wire [9:0] in_dat_wire64  = in_dat_wire[4489:4480] ;
    wire [9:0] in_dat_wire65  = in_dat_wire[4479:4470] ;
    wire [9:0] in_dat_wire66  = in_dat_wire[4469:4460] ;
    wire [9:0] in_dat_wire67  = in_dat_wire[4459:4450] ;
    wire [9:0] in_dat_wire68  = in_dat_wire[4449:4440] ;
    wire [9:0] in_dat_wire69  = in_dat_wire[4439:4430] ;
    wire [9:0] in_dat_wire70  = in_dat_wire[4429:4420] ;
    wire [9:0] in_dat_wire71  = in_dat_wire[4419:4410] ;
    wire [9:0] in_dat_wire72  = in_dat_wire[4409:4400] ;
    wire [9:0] in_dat_wire73  = in_dat_wire[4399:4390] ;
    wire [9:0] in_dat_wire74  = in_dat_wire[4389:4380] ;
    wire [9:0] in_dat_wire75  = in_dat_wire[4379:4370] ;
    wire [9:0] in_dat_wire76  = in_dat_wire[4369:4360] ;
    wire [9:0] in_dat_wire77  = in_dat_wire[4359:4350] ;
    wire [9:0] in_dat_wire78  = in_dat_wire[4349:4340] ;
    wire [9:0] in_dat_wire79  = in_dat_wire[4339:4330] ;
    wire [9:0] in_dat_wire80  = in_dat_wire[4329:4320] ;
    wire [9:0] in_dat_wire81  = in_dat_wire[4319:4310] ;
    wire [9:0] in_dat_wire82  = in_dat_wire[4309:4300] ;
    wire [9:0] in_dat_wire83  = in_dat_wire[4299:4290] ;
    wire [9:0] in_dat_wire84  = in_dat_wire[4289:4280] ;
    wire [9:0] in_dat_wire85  = in_dat_wire[4279:4270] ;
    wire [9:0] in_dat_wire86  = in_dat_wire[4269:4260] ;
    wire [9:0] in_dat_wire87  = in_dat_wire[4259:4250] ;
    wire [9:0] in_dat_wire88  = in_dat_wire[4249:4240] ;
    wire [9:0] in_dat_wire89  = in_dat_wire[4239:4230] ;
    wire [9:0] in_dat_wire90  = in_dat_wire[4229:4220] ;
    wire [9:0] in_dat_wire91  = in_dat_wire[4219:4210] ;
    wire [9:0] in_dat_wire92  = in_dat_wire[4209:4200] ;
    wire [9:0] in_dat_wire93  = in_dat_wire[4199:4190] ;
    wire [9:0] in_dat_wire94  = in_dat_wire[4189:4180] ;
    wire [9:0] in_dat_wire95  = in_dat_wire[4179:4170] ;
    wire [9:0] in_dat_wire96  = in_dat_wire[4169:4160] ;
    wire [9:0] in_dat_wire97  = in_dat_wire[4159:4150] ;
    wire [9:0] in_dat_wire98  = in_dat_wire[4149:4140] ;
    wire [9:0] in_dat_wire99  = in_dat_wire[4139:4130] ;
    wire [9:0] in_dat_wire100 = in_dat_wire[4129:4120] ;
    wire [9:0] in_dat_wire101 = in_dat_wire[4119:4110] ;
    wire [9:0] in_dat_wire102 = in_dat_wire[4109:4100] ;
    wire [9:0] in_dat_wire103 = in_dat_wire[4099:4090] ;
    wire [9:0] in_dat_wire104 = in_dat_wire[4089:4080] ;
    wire [9:0] in_dat_wire105 = in_dat_wire[4079:4070] ;
    wire [9:0] in_dat_wire106 = in_dat_wire[4069:4060] ;
    wire [9:0] in_dat_wire107 = in_dat_wire[4059:4050] ;
    wire [9:0] in_dat_wire108 = in_dat_wire[4049:4040] ;
    wire [9:0] in_dat_wire109 = in_dat_wire[4039:4030] ;
    wire [9:0] in_dat_wire110 = in_dat_wire[4029:4020] ;
    wire [9:0] in_dat_wire111 = in_dat_wire[4019:4010] ;
    wire [9:0] in_dat_wire112 = in_dat_wire[4009:4000] ;
    wire [9:0] in_dat_wire113 = in_dat_wire[3999:3990] ;
    wire [9:0] in_dat_wire114 = in_dat_wire[3989:3980] ;
    wire [9:0] in_dat_wire115 = in_dat_wire[3979:3970] ;
    wire [9:0] in_dat_wire116 = in_dat_wire[3969:3960] ;
    wire [9:0] in_dat_wire117 = in_dat_wire[3959:3950] ;
    wire [9:0] in_dat_wire118 = in_dat_wire[3949:3940] ;
    wire [9:0] in_dat_wire119 = in_dat_wire[3939:3930] ;
    wire [9:0] in_dat_wire120 = in_dat_wire[3929:3920] ;
    wire [9:0] in_dat_wire121 = in_dat_wire[3919:3910] ;
    wire [9:0] in_dat_wire122 = in_dat_wire[3909:3900] ;
    wire [9:0] in_dat_wire123 = in_dat_wire[3899:3890] ;
    wire [9:0] in_dat_wire124 = in_dat_wire[3889:3880] ;
    wire [9:0] in_dat_wire125 = in_dat_wire[3879:3870] ;
    wire [9:0] in_dat_wire126 = in_dat_wire[3869:3860] ;
    wire [9:0] in_dat_wire127 = in_dat_wire[3859:3850] ;
    wire [9:0] in_dat_wire128 = in_dat_wire[3849:3840] ;
    wire [9:0] in_dat_wire129 = in_dat_wire[3839:3830] ;
    wire [9:0] in_dat_wire130 = in_dat_wire[3829:3820] ;
    wire [9:0] in_dat_wire131 = in_dat_wire[3819:3810] ;
    wire [9:0] in_dat_wire132 = in_dat_wire[3809:3800] ;
    wire [9:0] in_dat_wire133 = in_dat_wire[3799:3790] ;
    wire [9:0] in_dat_wire134 = in_dat_wire[3789:3780] ;
    wire [9:0] in_dat_wire135 = in_dat_wire[3779:3770] ;
    wire [9:0] in_dat_wire136 = in_dat_wire[3769:3760] ;
    wire [9:0] in_dat_wire137 = in_dat_wire[3759:3750] ;
    wire [9:0] in_dat_wire138 = in_dat_wire[3749:3740] ;
    wire [9:0] in_dat_wire139 = in_dat_wire[3739:3730] ;
    wire [9:0] in_dat_wire140 = in_dat_wire[3729:3720] ;
    wire [9:0] in_dat_wire141 = in_dat_wire[3719:3710] ;
    wire [9:0] in_dat_wire142 = in_dat_wire[3709:3700] ;
    wire [9:0] in_dat_wire143 = in_dat_wire[3699:3690] ;
    wire [9:0] in_dat_wire144 = in_dat_wire[3689:3680] ;
    wire [9:0] in_dat_wire145 = in_dat_wire[3679:3670] ;
    wire [9:0] in_dat_wire146 = in_dat_wire[3669:3660] ;
    wire [9:0] in_dat_wire147 = in_dat_wire[3659:3650] ;
    wire [9:0] in_dat_wire148 = in_dat_wire[3649:3640] ;
    wire [9:0] in_dat_wire149 = in_dat_wire[3639:3630] ;
    wire [9:0] in_dat_wire150 = in_dat_wire[3629:3620] ;
    wire [9:0] in_dat_wire151 = in_dat_wire[3619:3610] ;
    wire [9:0] in_dat_wire152 = in_dat_wire[3609:3600] ;
    wire [9:0] in_dat_wire153 = in_dat_wire[3599:3590] ;
    wire [9:0] in_dat_wire154 = in_dat_wire[3589:3580] ;
    wire [9:0] in_dat_wire155 = in_dat_wire[3579:3570] ;
    wire [9:0] in_dat_wire156 = in_dat_wire[3569:3560] ;
    wire [9:0] in_dat_wire157 = in_dat_wire[3559:3550] ;
    wire [9:0] in_dat_wire158 = in_dat_wire[3549:3540] ;
    wire [9:0] in_dat_wire159 = in_dat_wire[3539:3530] ;
    wire [9:0] in_dat_wire160 = in_dat_wire[3529:3520] ;
    wire [9:0] in_dat_wire161 = in_dat_wire[3519:3510] ;
    wire [9:0] in_dat_wire162 = in_dat_wire[3509:3500] ;
    wire [9:0] in_dat_wire163 = in_dat_wire[3499:3490] ;
    wire [9:0] in_dat_wire164 = in_dat_wire[3489:3480] ;
    wire [9:0] in_dat_wire165 = in_dat_wire[3479:3470] ;
    wire [9:0] in_dat_wire166 = in_dat_wire[3469:3460] ;
    wire [9:0] in_dat_wire167 = in_dat_wire[3459:3450] ;
    wire [9:0] in_dat_wire168 = in_dat_wire[3449:3440] ;
    wire [9:0] in_dat_wire169 = in_dat_wire[3439:3430] ;
    wire [9:0] in_dat_wire170 = in_dat_wire[3429:3420] ;
    wire [9:0] in_dat_wire171 = in_dat_wire[3419:3410] ;
    wire [9:0] in_dat_wire172 = in_dat_wire[3409:3400] ;
    wire [9:0] in_dat_wire173 = in_dat_wire[3399:3390] ;
    wire [9:0] in_dat_wire174 = in_dat_wire[3389:3380] ;
    wire [9:0] in_dat_wire175 = in_dat_wire[3379:3370] ;
    wire [9:0] in_dat_wire176 = in_dat_wire[3369:3360] ;
    wire [9:0] in_dat_wire177 = in_dat_wire[3359:3350] ;
    wire [9:0] in_dat_wire178 = in_dat_wire[3349:3340] ;
    wire [9:0] in_dat_wire179 = in_dat_wire[3339:3330] ;
    wire [9:0] in_dat_wire180 = in_dat_wire[3329:3320] ;
    wire [9:0] in_dat_wire181 = in_dat_wire[3319:3310] ;
    wire [9:0] in_dat_wire182 = in_dat_wire[3309:3300] ;
    wire [9:0] in_dat_wire183 = in_dat_wire[3299:3290] ;
    wire [9:0] in_dat_wire184 = in_dat_wire[3289:3280] ;
    wire [9:0] in_dat_wire185 = in_dat_wire[3279:3270] ;
    wire [9:0] in_dat_wire186 = in_dat_wire[3269:3260] ;
    wire [9:0] in_dat_wire187 = in_dat_wire[3259:3250] ;
    wire [9:0] in_dat_wire188 = in_dat_wire[3249:3240] ;
    wire [9:0] in_dat_wire189 = in_dat_wire[3239:3230] ;
    wire [9:0] in_dat_wire190 = in_dat_wire[3229:3220] ;
    wire [9:0] in_dat_wire191 = in_dat_wire[3219:3210] ;
    wire [9:0] in_dat_wire192 = in_dat_wire[3209:3200] ;
    wire [9:0] in_dat_wire193 = in_dat_wire[3199:3190] ;
    wire [9:0] in_dat_wire194 = in_dat_wire[3189:3180] ;
    wire [9:0] in_dat_wire195 = in_dat_wire[3179:3170] ;
    wire [9:0] in_dat_wire196 = in_dat_wire[3169:3160] ;
    wire [9:0] in_dat_wire197 = in_dat_wire[3159:3150] ;
    wire [9:0] in_dat_wire198 = in_dat_wire[3149:3140] ;
    wire [9:0] in_dat_wire199 = in_dat_wire[3139:3130] ;
    wire [9:0] in_dat_wire200 = in_dat_wire[3129:3120] ;
    wire [9:0] in_dat_wire201 = in_dat_wire[3119:3110] ;
    wire [9:0] in_dat_wire202 = in_dat_wire[3109:3100] ;
    wire [9:0] in_dat_wire203 = in_dat_wire[3099:3090] ;
    wire [9:0] in_dat_wire204 = in_dat_wire[3089:3080] ;
    wire [9:0] in_dat_wire205 = in_dat_wire[3079:3070] ;
    wire [9:0] in_dat_wire206 = in_dat_wire[3069:3060] ;
    wire [9:0] in_dat_wire207 = in_dat_wire[3059:3050] ;
    wire [9:0] in_dat_wire208 = in_dat_wire[3049:3040] ;
    wire [9:0] in_dat_wire209 = in_dat_wire[3039:3030] ;
    wire [9:0] in_dat_wire210 = in_dat_wire[3029:3020] ;
    wire [9:0] in_dat_wire211 = in_dat_wire[3019:3010] ;
    wire [9:0] in_dat_wire212 = in_dat_wire[3009:3000] ;
    wire [9:0] in_dat_wire213 = in_dat_wire[2999:2990] ;
    wire [9:0] in_dat_wire214 = in_dat_wire[2989:2980] ;
    wire [9:0] in_dat_wire215 = in_dat_wire[2979:2970] ;
    wire [9:0] in_dat_wire216 = in_dat_wire[2969:2960] ;
    wire [9:0] in_dat_wire217 = in_dat_wire[2959:2950] ;
    wire [9:0] in_dat_wire218 = in_dat_wire[2949:2940] ;
    wire [9:0] in_dat_wire219 = in_dat_wire[2939:2930] ;
    wire [9:0] in_dat_wire220 = in_dat_wire[2929:2920] ;
    wire [9:0] in_dat_wire221 = in_dat_wire[2919:2910] ;
    wire [9:0] in_dat_wire222 = in_dat_wire[2909:2900] ;
    wire [9:0] in_dat_wire223 = in_dat_wire[2899:2890] ;
    wire [9:0] in_dat_wire224 = in_dat_wire[2889:2880] ;
    wire [9:0] in_dat_wire225 = in_dat_wire[2879:2870] ;
    wire [9:0] in_dat_wire226 = in_dat_wire[2869:2860] ;
    wire [9:0] in_dat_wire227 = in_dat_wire[2859:2850] ;
    wire [9:0] in_dat_wire228 = in_dat_wire[2849:2840] ;
    wire [9:0] in_dat_wire229 = in_dat_wire[2839:2830] ;
    wire [9:0] in_dat_wire230 = in_dat_wire[2829:2820] ;
    wire [9:0] in_dat_wire231 = in_dat_wire[2819:2810] ;
    wire [9:0] in_dat_wire232 = in_dat_wire[2809:2800] ;
    wire [9:0] in_dat_wire233 = in_dat_wire[2799:2790] ;
    wire [9:0] in_dat_wire234 = in_dat_wire[2789:2780] ;
    wire [9:0] in_dat_wire235 = in_dat_wire[2779:2770] ;
    wire [9:0] in_dat_wire236 = in_dat_wire[2769:2760] ;
    wire [9:0] in_dat_wire237 = in_dat_wire[2759:2750] ;
    wire [9:0] in_dat_wire238 = in_dat_wire[2749:2740] ;
    wire [9:0] in_dat_wire239 = in_dat_wire[2739:2730] ;
    wire [9:0] in_dat_wire240 = in_dat_wire[2729:2720] ;
    wire [9:0] in_dat_wire241 = in_dat_wire[2719:2710] ;
    wire [9:0] in_dat_wire242 = in_dat_wire[2709:2700] ;
    wire [9:0] in_dat_wire243 = in_dat_wire[2699:2690] ;
    wire [9:0] in_dat_wire244 = in_dat_wire[2689:2680] ;
    wire [9:0] in_dat_wire245 = in_dat_wire[2679:2670] ;
    wire [9:0] in_dat_wire246 = in_dat_wire[2669:2660] ;
    wire [9:0] in_dat_wire247 = in_dat_wire[2659:2650] ;
    wire [9:0] in_dat_wire248 = in_dat_wire[2649:2640] ;
    wire [9:0] in_dat_wire249 = in_dat_wire[2639:2630] ;
    wire [9:0] in_dat_wire250 = in_dat_wire[2629:2620] ;
    wire [9:0] in_dat_wire251 = in_dat_wire[2619:2610] ;
    wire [9:0] in_dat_wire252 = in_dat_wire[2609:2600] ;
    wire [9:0] in_dat_wire253 = in_dat_wire[2599:2590] ;
    wire [9:0] in_dat_wire254 = in_dat_wire[2589:2580] ;
    wire [9:0] in_dat_wire255 = in_dat_wire[2579:2570] ;
    wire [9:0] in_dat_wire256 = in_dat_wire[2569:2560] ;
    wire [9:0] in_dat_wire257 = in_dat_wire[2559:2550] ;
    wire [9:0] in_dat_wire258 = in_dat_wire[2549:2540] ;
    wire [9:0] in_dat_wire259 = in_dat_wire[2539:2530] ;
    wire [9:0] in_dat_wire260 = in_dat_wire[2529:2520] ;
    wire [9:0] in_dat_wire261 = in_dat_wire[2519:2510] ;
    wire [9:0] in_dat_wire262 = in_dat_wire[2509:2500] ;
    wire [9:0] in_dat_wire263 = in_dat_wire[2499:2490] ;
    wire [9:0] in_dat_wire264 = in_dat_wire[2489:2480] ;
    wire [9:0] in_dat_wire265 = in_dat_wire[2479:2470] ;
    wire [9:0] in_dat_wire266 = in_dat_wire[2469:2460] ;
    wire [9:0] in_dat_wire267 = in_dat_wire[2459:2450] ;
    wire [9:0] in_dat_wire268 = in_dat_wire[2449:2440] ;
    wire [9:0] in_dat_wire269 = in_dat_wire[2439:2430] ;
    wire [9:0] in_dat_wire270 = in_dat_wire[2429:2420] ;
    wire [9:0] in_dat_wire271 = in_dat_wire[2419:2410] ;
    wire [9:0] in_dat_wire272 = in_dat_wire[2409:2400] ;
    wire [9:0] in_dat_wire273 = in_dat_wire[2399:2390] ;
    wire [9:0] in_dat_wire274 = in_dat_wire[2389:2380] ;
    wire [9:0] in_dat_wire275 = in_dat_wire[2379:2370] ;
    wire [9:0] in_dat_wire276 = in_dat_wire[2369:2360] ;
    wire [9:0] in_dat_wire277 = in_dat_wire[2359:2350] ;
    wire [9:0] in_dat_wire278 = in_dat_wire[2349:2340] ;
    wire [9:0] in_dat_wire279 = in_dat_wire[2339:2330] ;
    wire [9:0] in_dat_wire280 = in_dat_wire[2329:2320] ;
    wire [9:0] in_dat_wire281 = in_dat_wire[2319:2310] ;
    wire [9:0] in_dat_wire282 = in_dat_wire[2309:2300] ;
    wire [9:0] in_dat_wire283 = in_dat_wire[2299:2290] ;
    wire [9:0] in_dat_wire284 = in_dat_wire[2289:2280] ;
    wire [9:0] in_dat_wire285 = in_dat_wire[2279:2270] ;
    wire [9:0] in_dat_wire286 = in_dat_wire[2269:2260] ;
    wire [9:0] in_dat_wire287 = in_dat_wire[2259:2250] ;
    wire [9:0] in_dat_wire288 = in_dat_wire[2249:2240] ;
    wire [9:0] in_dat_wire289 = in_dat_wire[2239:2230] ;
    wire [9:0] in_dat_wire290 = in_dat_wire[2229:2220] ;
    wire [9:0] in_dat_wire291 = in_dat_wire[2219:2210] ;
    wire [9:0] in_dat_wire292 = in_dat_wire[2209:2200] ;
    wire [9:0] in_dat_wire293 = in_dat_wire[2199:2190] ;
    wire [9:0] in_dat_wire294 = in_dat_wire[2189:2180] ;
    wire [9:0] in_dat_wire295 = in_dat_wire[2179:2170] ;
    wire [9:0] in_dat_wire296 = in_dat_wire[2169:2160] ;
    wire [9:0] in_dat_wire297 = in_dat_wire[2159:2150] ;
    wire [9:0] in_dat_wire298 = in_dat_wire[2149:2140] ;
    wire [9:0] in_dat_wire299 = in_dat_wire[2139:2130] ;
    wire [9:0] in_dat_wire300 = in_dat_wire[2129:2120] ;
    wire [9:0] in_dat_wire301 = in_dat_wire[2119:2110] ;
    wire [9:0] in_dat_wire302 = in_dat_wire[2109:2100] ;
    wire [9:0] in_dat_wire303 = in_dat_wire[2099:2090] ;
    wire [9:0] in_dat_wire304 = in_dat_wire[2089:2080] ;
    wire [9:0] in_dat_wire305 = in_dat_wire[2079:2070] ;
    wire [9:0] in_dat_wire306 = in_dat_wire[2069:2060] ;
    wire [9:0] in_dat_wire307 = in_dat_wire[2059:2050] ;
    wire [9:0] in_dat_wire308 = in_dat_wire[2049:2040] ;
    wire [9:0] in_dat_wire309 = in_dat_wire[2039:2030] ;
    wire [9:0] in_dat_wire310 = in_dat_wire[2029:2020] ;
    wire [9:0] in_dat_wire311 = in_dat_wire[2019:2010] ;
    wire [9:0] in_dat_wire312 = in_dat_wire[2009:2000] ;
    wire [9:0] in_dat_wire313 = in_dat_wire[1999:1990] ;
    wire [9:0] in_dat_wire314 = in_dat_wire[1989:1980] ;
    wire [9:0] in_dat_wire315 = in_dat_wire[1979:1970] ;
    wire [9:0] in_dat_wire316 = in_dat_wire[1969:1960] ;
    wire [9:0] in_dat_wire317 = in_dat_wire[1959:1950] ;
    wire [9:0] in_dat_wire318 = in_dat_wire[1949:1940] ;
    wire [9:0] in_dat_wire319 = in_dat_wire[1939:1930] ;
    wire [9:0] in_dat_wire320 = in_dat_wire[1929:1920] ;
    wire [9:0] in_dat_wire321 = in_dat_wire[1919:1910] ;
    wire [9:0] in_dat_wire322 = in_dat_wire[1909:1900] ;
    wire [9:0] in_dat_wire323 = in_dat_wire[1899:1890] ;
    wire [9:0] in_dat_wire324 = in_dat_wire[1889:1880] ;
    wire [9:0] in_dat_wire325 = in_dat_wire[1879:1870] ;
    wire [9:0] in_dat_wire326 = in_dat_wire[1869:1860] ;
    wire [9:0] in_dat_wire327 = in_dat_wire[1859:1850] ;
    wire [9:0] in_dat_wire328 = in_dat_wire[1849:1840] ;
    wire [9:0] in_dat_wire329 = in_dat_wire[1839:1830] ;
    wire [9:0] in_dat_wire330 = in_dat_wire[1829:1820] ;
    wire [9:0] in_dat_wire331 = in_dat_wire[1819:1810] ;
    wire [9:0] in_dat_wire332 = in_dat_wire[1809:1800] ;
    wire [9:0] in_dat_wire333 = in_dat_wire[1799:1790] ;
    wire [9:0] in_dat_wire334 = in_dat_wire[1789:1780] ;
    wire [9:0] in_dat_wire335 = in_dat_wire[1779:1770] ;
    wire [9:0] in_dat_wire336 = in_dat_wire[1769:1760] ;
    wire [9:0] in_dat_wire337 = in_dat_wire[1759:1750] ;
    wire [9:0] in_dat_wire338 = in_dat_wire[1749:1740] ;
    wire [9:0] in_dat_wire339 = in_dat_wire[1739:1730] ;
    wire [9:0] in_dat_wire340 = in_dat_wire[1729:1720] ;
    wire [9:0] in_dat_wire341 = in_dat_wire[1719:1710] ;
    wire [9:0] in_dat_wire342 = in_dat_wire[1709:1700] ;
    wire [9:0] in_dat_wire343 = in_dat_wire[1699:1690] ;
    wire [9:0] in_dat_wire344 = in_dat_wire[1689:1680] ;
    wire [9:0] in_dat_wire345 = in_dat_wire[1679:1670] ;
    wire [9:0] in_dat_wire346 = in_dat_wire[1669:1660] ;
    wire [9:0] in_dat_wire347 = in_dat_wire[1659:1650] ;
    wire [9:0] in_dat_wire348 = in_dat_wire[1649:1640] ;
    wire [9:0] in_dat_wire349 = in_dat_wire[1639:1630] ;
    wire [9:0] in_dat_wire350 = in_dat_wire[1629:1620] ;
    wire [9:0] in_dat_wire351 = in_dat_wire[1619:1610] ;
    wire [9:0] in_dat_wire352 = in_dat_wire[1609:1600] ;
    wire [9:0] in_dat_wire353 = in_dat_wire[1599:1590] ;
    wire [9:0] in_dat_wire354 = in_dat_wire[1589:1580] ;
    wire [9:0] in_dat_wire355 = in_dat_wire[1579:1570] ;
    wire [9:0] in_dat_wire356 = in_dat_wire[1569:1560] ;
    wire [9:0] in_dat_wire357 = in_dat_wire[1559:1550] ;
    wire [9:0] in_dat_wire358 = in_dat_wire[1549:1540] ;
    wire [9:0] in_dat_wire359 = in_dat_wire[1539:1530] ;
    wire [9:0] in_dat_wire360 = in_dat_wire[1529:1520] ;
    wire [9:0] in_dat_wire361 = in_dat_wire[1519:1510] ;
    wire [9:0] in_dat_wire362 = in_dat_wire[1509:1500] ;
    wire [9:0] in_dat_wire363 = in_dat_wire[1499:1490] ;
    wire [9:0] in_dat_wire364 = in_dat_wire[1489:1480] ;
    wire [9:0] in_dat_wire365 = in_dat_wire[1479:1470] ;
    wire [9:0] in_dat_wire366 = in_dat_wire[1469:1460] ;
    wire [9:0] in_dat_wire367 = in_dat_wire[1459:1450] ;
    wire [9:0] in_dat_wire368 = in_dat_wire[1449:1440] ;
    wire [9:0] in_dat_wire369 = in_dat_wire[1439:1430] ;
    wire [9:0] in_dat_wire370 = in_dat_wire[1429:1420] ;
    wire [9:0] in_dat_wire371 = in_dat_wire[1419:1410] ;
    wire [9:0] in_dat_wire372 = in_dat_wire[1409:1400] ;
    wire [9:0] in_dat_wire373 = in_dat_wire[1399:1390] ;
    wire [9:0] in_dat_wire374 = in_dat_wire[1389:1380] ;
    wire [9:0] in_dat_wire375 = in_dat_wire[1379:1370] ;
    wire [9:0] in_dat_wire376 = in_dat_wire[1369:1360] ;
    wire [9:0] in_dat_wire377 = in_dat_wire[1359:1350] ;
    wire [9:0] in_dat_wire378 = in_dat_wire[1349:1340] ;
    wire [9:0] in_dat_wire379 = in_dat_wire[1339:1330] ;
    wire [9:0] in_dat_wire380 = in_dat_wire[1329:1320] ;
    wire [9:0] in_dat_wire381 = in_dat_wire[1319:1310] ;
    wire [9:0] in_dat_wire382 = in_dat_wire[1309:1300] ;
    wire [9:0] in_dat_wire383 = in_dat_wire[1299:1290] ;
    wire [9:0] in_dat_wire384 = in_dat_wire[1289:1280] ;
    wire [9:0] in_dat_wire385 = in_dat_wire[1279:1270] ;
    wire [9:0] in_dat_wire386 = in_dat_wire[1269:1260] ;
    wire [9:0] in_dat_wire387 = in_dat_wire[1259:1250] ;
    wire [9:0] in_dat_wire388 = in_dat_wire[1249:1240] ;
    wire [9:0] in_dat_wire389 = in_dat_wire[1239:1230] ;
    wire [9:0] in_dat_wire390 = in_dat_wire[1229:1220] ;
    wire [9:0] in_dat_wire391 = in_dat_wire[1219:1210] ;
    wire [9:0] in_dat_wire392 = in_dat_wire[1209:1200] ;
    wire [9:0] in_dat_wire393 = in_dat_wire[1199:1190] ;
    wire [9:0] in_dat_wire394 = in_dat_wire[1189:1180] ;
    wire [9:0] in_dat_wire395 = in_dat_wire[1179:1170] ;
    wire [9:0] in_dat_wire396 = in_dat_wire[1169:1160] ;
    wire [9:0] in_dat_wire397 = in_dat_wire[1159:1150] ;
    wire [9:0] in_dat_wire398 = in_dat_wire[1149:1140] ;
    wire [9:0] in_dat_wire399 = in_dat_wire[1139:1130] ;
    wire [9:0] in_dat_wire400 = in_dat_wire[1129:1120] ;
    wire [9:0] in_dat_wire401 = in_dat_wire[1119:1110] ;
    wire [9:0] in_dat_wire402 = in_dat_wire[1109:1100] ;
    wire [9:0] in_dat_wire403 = in_dat_wire[1099:1090] ;
    wire [9:0] in_dat_wire404 = in_dat_wire[1089:1080] ;
    wire [9:0] in_dat_wire405 = in_dat_wire[1079:1070] ;
    wire [9:0] in_dat_wire406 = in_dat_wire[1069:1060] ;
    wire [9:0] in_dat_wire407 = in_dat_wire[1059:1050] ;
    wire [9:0] in_dat_wire408 = in_dat_wire[1049:1040] ;
    wire [9:0] in_dat_wire409 = in_dat_wire[1039:1030] ;
    wire [9:0] in_dat_wire410 = in_dat_wire[1029:1020] ;
    wire [9:0] in_dat_wire411 = in_dat_wire[1019:1010] ;
    wire [9:0] in_dat_wire412 = in_dat_wire[1009:1000] ;
    wire [9:0] in_dat_wire413 = in_dat_wire[999:990] ;
    wire [9:0] in_dat_wire414 = in_dat_wire[989:980] ;
    wire [9:0] in_dat_wire415 = in_dat_wire[979:970] ;
    wire [9:0] in_dat_wire416 = in_dat_wire[969:960] ;
    wire [9:0] in_dat_wire417 = in_dat_wire[959:950] ;
    wire [9:0] in_dat_wire418 = in_dat_wire[949:940] ;
    wire [9:0] in_dat_wire419 = in_dat_wire[939:930] ;
    wire [9:0] in_dat_wire420 = in_dat_wire[929:920] ;
    wire [9:0] in_dat_wire421 = in_dat_wire[919:910] ;
    wire [9:0] in_dat_wire422 = in_dat_wire[909:900] ;
    wire [9:0] in_dat_wire423 = in_dat_wire[899:890] ;
    wire [9:0] in_dat_wire424 = in_dat_wire[889:880] ;
    wire [9:0] in_dat_wire425 = in_dat_wire[879:870] ;
    wire [9:0] in_dat_wire426 = in_dat_wire[869:860] ;
    wire [9:0] in_dat_wire427 = in_dat_wire[859:850] ;
    wire [9:0] in_dat_wire428 = in_dat_wire[849:840] ;
    wire [9:0] in_dat_wire429 = in_dat_wire[839:830] ;
    wire [9:0] in_dat_wire430 = in_dat_wire[829:820] ;
    wire [9:0] in_dat_wire431 = in_dat_wire[819:810] ;
    wire [9:0] in_dat_wire432 = in_dat_wire[809:800] ;
    wire [9:0] in_dat_wire433 = in_dat_wire[799:790] ;
    wire [9:0] in_dat_wire434 = in_dat_wire[789:780] ;
    wire [9:0] in_dat_wire435 = in_dat_wire[779:770] ;
    wire [9:0] in_dat_wire436 = in_dat_wire[769:760] ;
    wire [9:0] in_dat_wire437 = in_dat_wire[759:750] ;
    wire [9:0] in_dat_wire438 = in_dat_wire[749:740] ;
    wire [9:0] in_dat_wire439 = in_dat_wire[739:730] ;
    wire [9:0] in_dat_wire440 = in_dat_wire[729:720] ;
    wire [9:0] in_dat_wire441 = in_dat_wire[719:710] ;
    wire [9:0] in_dat_wire442 = in_dat_wire[709:700] ;
    wire [9:0] in_dat_wire443 = in_dat_wire[699:690] ;
    wire [9:0] in_dat_wire444 = in_dat_wire[689:680] ;
    wire [9:0] in_dat_wire445 = in_dat_wire[679:670] ;
    wire [9:0] in_dat_wire446 = in_dat_wire[669:660] ;
    wire [9:0] in_dat_wire447 = in_dat_wire[659:650] ;
    wire [9:0] in_dat_wire448 = in_dat_wire[649:640] ;
    wire [9:0] in_dat_wire449 = in_dat_wire[639:630] ;
    wire [9:0] in_dat_wire450 = in_dat_wire[629:620] ;
    wire [9:0] in_dat_wire451 = in_dat_wire[619:610] ;
    wire [9:0] in_dat_wire452 = in_dat_wire[609:600] ;
    wire [9:0] in_dat_wire453 = in_dat_wire[599:590] ;
    wire [9:0] in_dat_wire454 = in_dat_wire[589:580] ;
    wire [9:0] in_dat_wire455 = in_dat_wire[579:570] ;
    wire [9:0] in_dat_wire456 = in_dat_wire[569:560] ;
    wire [9:0] in_dat_wire457 = in_dat_wire[559:550] ;
    wire [9:0] in_dat_wire458 = in_dat_wire[549:540] ;
    wire [9:0] in_dat_wire459 = in_dat_wire[539:530] ;
    wire [9:0] in_dat_wire460 = in_dat_wire[529:520] ;
    wire [9:0] in_dat_wire461 = in_dat_wire[519:510] ;
    wire [9:0] in_dat_wire462 = in_dat_wire[509:500] ;
    wire [9:0] in_dat_wire463 = in_dat_wire[499:490] ;
    wire [9:0] in_dat_wire464 = in_dat_wire[489:480] ;
    wire [9:0] in_dat_wire465 = in_dat_wire[479:470] ;
    wire [9:0] in_dat_wire466 = in_dat_wire[469:460] ;
    wire [9:0] in_dat_wire467 = in_dat_wire[459:450] ;
    wire [9:0] in_dat_wire468 = in_dat_wire[449:440] ;
    wire [9:0] in_dat_wire469 = in_dat_wire[439:430] ;
    wire [9:0] in_dat_wire470 = in_dat_wire[429:420] ;
    wire [9:0] in_dat_wire471 = in_dat_wire[419:410] ;
    wire [9:0] in_dat_wire472 = in_dat_wire[409:400] ;
    wire [9:0] in_dat_wire473 = in_dat_wire[399:390] ;
    wire [9:0] in_dat_wire474 = in_dat_wire[389:380] ;
    wire [9:0] in_dat_wire475 = in_dat_wire[379:370] ;
    wire [9:0] in_dat_wire476 = in_dat_wire[369:360] ;
    wire [9:0] in_dat_wire477 = in_dat_wire[359:350] ;
    wire [9:0] in_dat_wire478 = in_dat_wire[349:340] ;
    wire [9:0] in_dat_wire479 = in_dat_wire[339:330] ;
    wire [9:0] in_dat_wire480 = in_dat_wire[329:320] ;
    wire [9:0] in_dat_wire481 = in_dat_wire[319:310] ;
    wire [9:0] in_dat_wire482 = in_dat_wire[309:300] ;
    wire [9:0] in_dat_wire483 = in_dat_wire[299:290] ;
    wire [9:0] in_dat_wire484 = in_dat_wire[289:280] ;
    wire [9:0] in_dat_wire485 = in_dat_wire[279:270] ;
    wire [9:0] in_dat_wire486 = in_dat_wire[269:260] ;
    wire [9:0] in_dat_wire487 = in_dat_wire[259:250] ;
    wire [9:0] in_dat_wire488 = in_dat_wire[249:240] ;
    wire [9:0] in_dat_wire489 = in_dat_wire[239:230] ;
    wire [9:0] in_dat_wire490 = in_dat_wire[229:220] ;
    wire [9:0] in_dat_wire491 = in_dat_wire[219:210] ;
    wire [9:0] in_dat_wire492 = in_dat_wire[209:200] ;
    wire [9:0] in_dat_wire493 = in_dat_wire[199:190] ;
    wire [9:0] in_dat_wire494 = in_dat_wire[189:180] ;
    wire [9:0] in_dat_wire495 = in_dat_wire[179:170] ;
    wire [9:0] in_dat_wire496 = in_dat_wire[169:160] ;
    wire [9:0] in_dat_wire497 = in_dat_wire[159:150] ;
    wire [9:0] in_dat_wire498 = in_dat_wire[149:140] ;
    wire [9:0] in_dat_wire499 = in_dat_wire[139:130] ;
    wire [9:0] in_dat_wire500 = in_dat_wire[129:120] ;
    wire [9:0] in_dat_wire501 = in_dat_wire[119:110] ;
    wire [9:0] in_dat_wire502 = in_dat_wire[109:100] ;
    wire [9:0] in_dat_wire503 = in_dat_wire[99:90] ;
    wire [9:0] in_dat_wire504 = in_dat_wire[89:80] ;
    wire [9:0] in_dat_wire505 = in_dat_wire[79:70] ;
    wire [9:0] in_dat_wire506 = in_dat_wire[69:60] ;
    wire [9:0] in_dat_wire507 = in_dat_wire[59:50] ;
    wire [9:0] in_dat_wire508 = in_dat_wire[49:40] ;
    wire [9:0] in_dat_wire509 = in_dat_wire[39:30] ;
    wire [9:0] in_dat_wire510 = in_dat_wire[29:20] ;
    wire [9:0] in_dat_wire511 = in_dat_wire[19:10] ;
    wire [9:0] in_dat_wire512 = in_dat_wire[9:0] ;

    wire [9:0] coe_dat_wire01  = coe_dat_wire[5119:5110] ;
    wire [9:0] coe_dat_wire02  = coe_dat_wire[5109:5100] ;
    wire [9:0] coe_dat_wire03  = coe_dat_wire[5099:5090] ;
    wire [9:0] coe_dat_wire04  = coe_dat_wire[5089:5080] ;
    wire [9:0] coe_dat_wire05  = coe_dat_wire[5079:5070] ;
    wire [9:0] coe_dat_wire06  = coe_dat_wire[5069:5060] ;
    wire [9:0] coe_dat_wire07  = coe_dat_wire[5059:5050] ;
    wire [9:0] coe_dat_wire08  = coe_dat_wire[5049:5040] ;
    wire [9:0] coe_dat_wire09  = coe_dat_wire[5039:5030] ;
    wire [9:0] coe_dat_wire10  = coe_dat_wire[5029:5020] ;
    wire [9:0] coe_dat_wire11  = coe_dat_wire[5019:5010] ;
    wire [9:0] coe_dat_wire12  = coe_dat_wire[5009:5000] ;
    wire [9:0] coe_dat_wire13  = coe_dat_wire[4999:4990] ;
    wire [9:0] coe_dat_wire14  = coe_dat_wire[4989:4980] ;
    wire [9:0] coe_dat_wire15  = coe_dat_wire[4979:4970] ;
    wire [9:0] coe_dat_wire16  = coe_dat_wire[4969:4960] ;
    wire [9:0] coe_dat_wire17  = coe_dat_wire[4959:4950] ;
    wire [9:0] coe_dat_wire18  = coe_dat_wire[4949:4940] ;
    wire [9:0] coe_dat_wire19  = coe_dat_wire[4939:4930] ;
    wire [9:0] coe_dat_wire20  = coe_dat_wire[4929:4920] ;
    wire [9:0] coe_dat_wire21  = coe_dat_wire[4919:4910] ;
    wire [9:0] coe_dat_wire22  = coe_dat_wire[4909:4900] ;
    wire [9:0] coe_dat_wire23  = coe_dat_wire[4899:4890] ;
    wire [9:0] coe_dat_wire24  = coe_dat_wire[4889:4880] ;
    wire [9:0] coe_dat_wire25  = coe_dat_wire[4879:4870] ;
    wire [9:0] coe_dat_wire26  = coe_dat_wire[4869:4860] ;
    wire [9:0] coe_dat_wire27  = coe_dat_wire[4859:4850] ;
    wire [9:0] coe_dat_wire28  = coe_dat_wire[4849:4840] ;
    wire [9:0] coe_dat_wire29  = coe_dat_wire[4839:4830] ;
    wire [9:0] coe_dat_wire30  = coe_dat_wire[4829:4820] ;
    wire [9:0] coe_dat_wire31  = coe_dat_wire[4819:4810] ;
    wire [9:0] coe_dat_wire32  = coe_dat_wire[4809:4800] ;
    wire [9:0] coe_dat_wire33  = coe_dat_wire[4799:4790] ;
    wire [9:0] coe_dat_wire34  = coe_dat_wire[4789:4780] ;
    wire [9:0] coe_dat_wire35  = coe_dat_wire[4779:4770] ;
    wire [9:0] coe_dat_wire36  = coe_dat_wire[4769:4760] ;
    wire [9:0] coe_dat_wire37  = coe_dat_wire[4759:4750] ;
    wire [9:0] coe_dat_wire38  = coe_dat_wire[4749:4740] ;
    wire [9:0] coe_dat_wire39  = coe_dat_wire[4739:4730] ;
    wire [9:0] coe_dat_wire40  = coe_dat_wire[4729:4720] ;
    wire [9:0] coe_dat_wire41  = coe_dat_wire[4719:4710] ;
    wire [9:0] coe_dat_wire42  = coe_dat_wire[4709:4700] ;
    wire [9:0] coe_dat_wire43  = coe_dat_wire[4699:4690] ;
    wire [9:0] coe_dat_wire44  = coe_dat_wire[4689:4680] ;
    wire [9:0] coe_dat_wire45  = coe_dat_wire[4679:4670] ;
    wire [9:0] coe_dat_wire46  = coe_dat_wire[4669:4660] ;
    wire [9:0] coe_dat_wire47  = coe_dat_wire[4659:4650] ;
    wire [9:0] coe_dat_wire48  = coe_dat_wire[4649:4640] ;
    wire [9:0] coe_dat_wire49  = coe_dat_wire[4639:4630] ;
    wire [9:0] coe_dat_wire50  = coe_dat_wire[4629:4620] ;
    wire [9:0] coe_dat_wire51  = coe_dat_wire[4619:4610] ;
    wire [9:0] coe_dat_wire52  = coe_dat_wire[4609:4600] ;
    wire [9:0] coe_dat_wire53  = coe_dat_wire[4599:4590] ;
    wire [9:0] coe_dat_wire54  = coe_dat_wire[4589:4580] ;
    wire [9:0] coe_dat_wire55  = coe_dat_wire[4579:4570] ;
    wire [9:0] coe_dat_wire56  = coe_dat_wire[4569:4560] ;
    wire [9:0] coe_dat_wire57  = coe_dat_wire[4559:4550] ;
    wire [9:0] coe_dat_wire58  = coe_dat_wire[4549:4540] ;
    wire [9:0] coe_dat_wire59  = coe_dat_wire[4539:4530] ;
    wire [9:0] coe_dat_wire60  = coe_dat_wire[4529:4520] ;
    wire [9:0] coe_dat_wire61  = coe_dat_wire[4519:4510] ;
    wire [9:0] coe_dat_wire62  = coe_dat_wire[4509:4500] ;
    wire [9:0] coe_dat_wire63  = coe_dat_wire[4499:4490] ;
    wire [9:0] coe_dat_wire64  = coe_dat_wire[4489:4480] ;
    wire [9:0] coe_dat_wire65  = coe_dat_wire[4479:4470] ;
    wire [9:0] coe_dat_wire66  = coe_dat_wire[4469:4460] ;
    wire [9:0] coe_dat_wire67  = coe_dat_wire[4459:4450] ;
    wire [9:0] coe_dat_wire68  = coe_dat_wire[4449:4440] ;
    wire [9:0] coe_dat_wire69  = coe_dat_wire[4439:4430] ;
    wire [9:0] coe_dat_wire70  = coe_dat_wire[4429:4420] ;
    wire [9:0] coe_dat_wire71  = coe_dat_wire[4419:4410] ;
    wire [9:0] coe_dat_wire72  = coe_dat_wire[4409:4400] ;
    wire [9:0] coe_dat_wire73  = coe_dat_wire[4399:4390] ;
    wire [9:0] coe_dat_wire74  = coe_dat_wire[4389:4380] ;
    wire [9:0] coe_dat_wire75  = coe_dat_wire[4379:4370] ;
    wire [9:0] coe_dat_wire76  = coe_dat_wire[4369:4360] ;
    wire [9:0] coe_dat_wire77  = coe_dat_wire[4359:4350] ;
    wire [9:0] coe_dat_wire78  = coe_dat_wire[4349:4340] ;
    wire [9:0] coe_dat_wire79  = coe_dat_wire[4339:4330] ;
    wire [9:0] coe_dat_wire80  = coe_dat_wire[4329:4320] ;
    wire [9:0] coe_dat_wire81  = coe_dat_wire[4319:4310] ;
    wire [9:0] coe_dat_wire82  = coe_dat_wire[4309:4300] ;
    wire [9:0] coe_dat_wire83  = coe_dat_wire[4299:4290] ;
    wire [9:0] coe_dat_wire84  = coe_dat_wire[4289:4280] ;
    wire [9:0] coe_dat_wire85  = coe_dat_wire[4279:4270] ;
    wire [9:0] coe_dat_wire86  = coe_dat_wire[4269:4260] ;
    wire [9:0] coe_dat_wire87  = coe_dat_wire[4259:4250] ;
    wire [9:0] coe_dat_wire88  = coe_dat_wire[4249:4240] ;
    wire [9:0] coe_dat_wire89  = coe_dat_wire[4239:4230] ;
    wire [9:0] coe_dat_wire90  = coe_dat_wire[4229:4220] ;
    wire [9:0] coe_dat_wire91  = coe_dat_wire[4219:4210] ;
    wire [9:0] coe_dat_wire92  = coe_dat_wire[4209:4200] ;
    wire [9:0] coe_dat_wire93  = coe_dat_wire[4199:4190] ;
    wire [9:0] coe_dat_wire94  = coe_dat_wire[4189:4180] ;
    wire [9:0] coe_dat_wire95  = coe_dat_wire[4179:4170] ;
    wire [9:0] coe_dat_wire96  = coe_dat_wire[4169:4160] ;
    wire [9:0] coe_dat_wire97  = coe_dat_wire[4159:4150] ;
    wire [9:0] coe_dat_wire98  = coe_dat_wire[4149:4140] ;
    wire [9:0] coe_dat_wire99  = coe_dat_wire[4139:4130] ;
    wire [9:0] coe_dat_wire100 = coe_dat_wire[4129:4120] ;
    wire [9:0] coe_dat_wire101 = coe_dat_wire[4119:4110] ;
    wire [9:0] coe_dat_wire102 = coe_dat_wire[4109:4100] ;
    wire [9:0] coe_dat_wire103 = coe_dat_wire[4099:4090] ;
    wire [9:0] coe_dat_wire104 = coe_dat_wire[4089:4080] ;
    wire [9:0] coe_dat_wire105 = coe_dat_wire[4079:4070] ;
    wire [9:0] coe_dat_wire106 = coe_dat_wire[4069:4060] ;
    wire [9:0] coe_dat_wire107 = coe_dat_wire[4059:4050] ;
    wire [9:0] coe_dat_wire108 = coe_dat_wire[4049:4040] ;
    wire [9:0] coe_dat_wire109 = coe_dat_wire[4039:4030] ;
    wire [9:0] coe_dat_wire110 = coe_dat_wire[4029:4020] ;
    wire [9:0] coe_dat_wire111 = coe_dat_wire[4019:4010] ;
    wire [9:0] coe_dat_wire112 = coe_dat_wire[4009:4000] ;
    wire [9:0] coe_dat_wire113 = coe_dat_wire[3999:3990] ;
    wire [9:0] coe_dat_wire114 = coe_dat_wire[3989:3980] ;
    wire [9:0] coe_dat_wire115 = coe_dat_wire[3979:3970] ;
    wire [9:0] coe_dat_wire116 = coe_dat_wire[3969:3960] ;
    wire [9:0] coe_dat_wire117 = coe_dat_wire[3959:3950] ;
    wire [9:0] coe_dat_wire118 = coe_dat_wire[3949:3940] ;
    wire [9:0] coe_dat_wire119 = coe_dat_wire[3939:3930] ;
    wire [9:0] coe_dat_wire120 = coe_dat_wire[3929:3920] ;
    wire [9:0] coe_dat_wire121 = coe_dat_wire[3919:3910] ;
    wire [9:0] coe_dat_wire122 = coe_dat_wire[3909:3900] ;
    wire [9:0] coe_dat_wire123 = coe_dat_wire[3899:3890] ;
    wire [9:0] coe_dat_wire124 = coe_dat_wire[3889:3880] ;
    wire [9:0] coe_dat_wire125 = coe_dat_wire[3879:3870] ;
    wire [9:0] coe_dat_wire126 = coe_dat_wire[3869:3860] ;
    wire [9:0] coe_dat_wire127 = coe_dat_wire[3859:3850] ;
    wire [9:0] coe_dat_wire128 = coe_dat_wire[3849:3840] ;
    wire [9:0] coe_dat_wire129 = coe_dat_wire[3839:3830] ;
    wire [9:0] coe_dat_wire130 = coe_dat_wire[3829:3820] ;
    wire [9:0] coe_dat_wire131 = coe_dat_wire[3819:3810] ;
    wire [9:0] coe_dat_wire132 = coe_dat_wire[3809:3800] ;
    wire [9:0] coe_dat_wire133 = coe_dat_wire[3799:3790] ;
    wire [9:0] coe_dat_wire134 = coe_dat_wire[3789:3780] ;
    wire [9:0] coe_dat_wire135 = coe_dat_wire[3779:3770] ;
    wire [9:0] coe_dat_wire136 = coe_dat_wire[3769:3760] ;
    wire [9:0] coe_dat_wire137 = coe_dat_wire[3759:3750] ;
    wire [9:0] coe_dat_wire138 = coe_dat_wire[3749:3740] ;
    wire [9:0] coe_dat_wire139 = coe_dat_wire[3739:3730] ;
    wire [9:0] coe_dat_wire140 = coe_dat_wire[3729:3720] ;
    wire [9:0] coe_dat_wire141 = coe_dat_wire[3719:3710] ;
    wire [9:0] coe_dat_wire142 = coe_dat_wire[3709:3700] ;
    wire [9:0] coe_dat_wire143 = coe_dat_wire[3699:3690] ;
    wire [9:0] coe_dat_wire144 = coe_dat_wire[3689:3680] ;
    wire [9:0] coe_dat_wire145 = coe_dat_wire[3679:3670] ;
    wire [9:0] coe_dat_wire146 = coe_dat_wire[3669:3660] ;
    wire [9:0] coe_dat_wire147 = coe_dat_wire[3659:3650] ;
    wire [9:0] coe_dat_wire148 = coe_dat_wire[3649:3640] ;
    wire [9:0] coe_dat_wire149 = coe_dat_wire[3639:3630] ;
    wire [9:0] coe_dat_wire150 = coe_dat_wire[3629:3620] ;
    wire [9:0] coe_dat_wire151 = coe_dat_wire[3619:3610] ;
    wire [9:0] coe_dat_wire152 = coe_dat_wire[3609:3600] ;
    wire [9:0] coe_dat_wire153 = coe_dat_wire[3599:3590] ;
    wire [9:0] coe_dat_wire154 = coe_dat_wire[3589:3580] ;
    wire [9:0] coe_dat_wire155 = coe_dat_wire[3579:3570] ;
    wire [9:0] coe_dat_wire156 = coe_dat_wire[3569:3560] ;
    wire [9:0] coe_dat_wire157 = coe_dat_wire[3559:3550] ;
    wire [9:0] coe_dat_wire158 = coe_dat_wire[3549:3540] ;
    wire [9:0] coe_dat_wire159 = coe_dat_wire[3539:3530] ;
    wire [9:0] coe_dat_wire160 = coe_dat_wire[3529:3520] ;
    wire [9:0] coe_dat_wire161 = coe_dat_wire[3519:3510] ;
    wire [9:0] coe_dat_wire162 = coe_dat_wire[3509:3500] ;
    wire [9:0] coe_dat_wire163 = coe_dat_wire[3499:3490] ;
    wire [9:0] coe_dat_wire164 = coe_dat_wire[3489:3480] ;
    wire [9:0] coe_dat_wire165 = coe_dat_wire[3479:3470] ;
    wire [9:0] coe_dat_wire166 = coe_dat_wire[3469:3460] ;
    wire [9:0] coe_dat_wire167 = coe_dat_wire[3459:3450] ;
    wire [9:0] coe_dat_wire168 = coe_dat_wire[3449:3440] ;
    wire [9:0] coe_dat_wire169 = coe_dat_wire[3439:3430] ;
    wire [9:0] coe_dat_wire170 = coe_dat_wire[3429:3420] ;
    wire [9:0] coe_dat_wire171 = coe_dat_wire[3419:3410] ;
    wire [9:0] coe_dat_wire172 = coe_dat_wire[3409:3400] ;
    wire [9:0] coe_dat_wire173 = coe_dat_wire[3399:3390] ;
    wire [9:0] coe_dat_wire174 = coe_dat_wire[3389:3380] ;
    wire [9:0] coe_dat_wire175 = coe_dat_wire[3379:3370] ;
    wire [9:0] coe_dat_wire176 = coe_dat_wire[3369:3360] ;
    wire [9:0] coe_dat_wire177 = coe_dat_wire[3359:3350] ;
    wire [9:0] coe_dat_wire178 = coe_dat_wire[3349:3340] ;
    wire [9:0] coe_dat_wire179 = coe_dat_wire[3339:3330] ;
    wire [9:0] coe_dat_wire180 = coe_dat_wire[3329:3320] ;
    wire [9:0] coe_dat_wire181 = coe_dat_wire[3319:3310] ;
    wire [9:0] coe_dat_wire182 = coe_dat_wire[3309:3300] ;
    wire [9:0] coe_dat_wire183 = coe_dat_wire[3299:3290] ;
    wire [9:0] coe_dat_wire184 = coe_dat_wire[3289:3280] ;
    wire [9:0] coe_dat_wire185 = coe_dat_wire[3279:3270] ;
    wire [9:0] coe_dat_wire186 = coe_dat_wire[3269:3260] ;
    wire [9:0] coe_dat_wire187 = coe_dat_wire[3259:3250] ;
    wire [9:0] coe_dat_wire188 = coe_dat_wire[3249:3240] ;
    wire [9:0] coe_dat_wire189 = coe_dat_wire[3239:3230] ;
    wire [9:0] coe_dat_wire190 = coe_dat_wire[3229:3220] ;
    wire [9:0] coe_dat_wire191 = coe_dat_wire[3219:3210] ;
    wire [9:0] coe_dat_wire192 = coe_dat_wire[3209:3200] ;
    wire [9:0] coe_dat_wire193 = coe_dat_wire[3199:3190] ;
    wire [9:0] coe_dat_wire194 = coe_dat_wire[3189:3180] ;
    wire [9:0] coe_dat_wire195 = coe_dat_wire[3179:3170] ;
    wire [9:0] coe_dat_wire196 = coe_dat_wire[3169:3160] ;
    wire [9:0] coe_dat_wire197 = coe_dat_wire[3159:3150] ;
    wire [9:0] coe_dat_wire198 = coe_dat_wire[3149:3140] ;
    wire [9:0] coe_dat_wire199 = coe_dat_wire[3139:3130] ;
    wire [9:0] coe_dat_wire200 = coe_dat_wire[3129:3120] ;
    wire [9:0] coe_dat_wire201 = coe_dat_wire[3119:3110] ;
    wire [9:0] coe_dat_wire202 = coe_dat_wire[3109:3100] ;
    wire [9:0] coe_dat_wire203 = coe_dat_wire[3099:3090] ;
    wire [9:0] coe_dat_wire204 = coe_dat_wire[3089:3080] ;
    wire [9:0] coe_dat_wire205 = coe_dat_wire[3079:3070] ;
    wire [9:0] coe_dat_wire206 = coe_dat_wire[3069:3060] ;
    wire [9:0] coe_dat_wire207 = coe_dat_wire[3059:3050] ;
    wire [9:0] coe_dat_wire208 = coe_dat_wire[3049:3040] ;
    wire [9:0] coe_dat_wire209 = coe_dat_wire[3039:3030] ;
    wire [9:0] coe_dat_wire210 = coe_dat_wire[3029:3020] ;
    wire [9:0] coe_dat_wire211 = coe_dat_wire[3019:3010] ;
    wire [9:0] coe_dat_wire212 = coe_dat_wire[3009:3000] ;
    wire [9:0] coe_dat_wire213 = coe_dat_wire[2999:2990] ;
    wire [9:0] coe_dat_wire214 = coe_dat_wire[2989:2980] ;
    wire [9:0] coe_dat_wire215 = coe_dat_wire[2979:2970] ;
    wire [9:0] coe_dat_wire216 = coe_dat_wire[2969:2960] ;
    wire [9:0] coe_dat_wire217 = coe_dat_wire[2959:2950] ;
    wire [9:0] coe_dat_wire218 = coe_dat_wire[2949:2940] ;
    wire [9:0] coe_dat_wire219 = coe_dat_wire[2939:2930] ;
    wire [9:0] coe_dat_wire220 = coe_dat_wire[2929:2920] ;
    wire [9:0] coe_dat_wire221 = coe_dat_wire[2919:2910] ;
    wire [9:0] coe_dat_wire222 = coe_dat_wire[2909:2900] ;
    wire [9:0] coe_dat_wire223 = coe_dat_wire[2899:2890] ;
    wire [9:0] coe_dat_wire224 = coe_dat_wire[2889:2880] ;
    wire [9:0] coe_dat_wire225 = coe_dat_wire[2879:2870] ;
    wire [9:0] coe_dat_wire226 = coe_dat_wire[2869:2860] ;
    wire [9:0] coe_dat_wire227 = coe_dat_wire[2859:2850] ;
    wire [9:0] coe_dat_wire228 = coe_dat_wire[2849:2840] ;
    wire [9:0] coe_dat_wire229 = coe_dat_wire[2839:2830] ;
    wire [9:0] coe_dat_wire230 = coe_dat_wire[2829:2820] ;
    wire [9:0] coe_dat_wire231 = coe_dat_wire[2819:2810] ;
    wire [9:0] coe_dat_wire232 = coe_dat_wire[2809:2800] ;
    wire [9:0] coe_dat_wire233 = coe_dat_wire[2799:2790] ;
    wire [9:0] coe_dat_wire234 = coe_dat_wire[2789:2780] ;
    wire [9:0] coe_dat_wire235 = coe_dat_wire[2779:2770] ;
    wire [9:0] coe_dat_wire236 = coe_dat_wire[2769:2760] ;
    wire [9:0] coe_dat_wire237 = coe_dat_wire[2759:2750] ;
    wire [9:0] coe_dat_wire238 = coe_dat_wire[2749:2740] ;
    wire [9:0] coe_dat_wire239 = coe_dat_wire[2739:2730] ;
    wire [9:0] coe_dat_wire240 = coe_dat_wire[2729:2720] ;
    wire [9:0] coe_dat_wire241 = coe_dat_wire[2719:2710] ;
    wire [9:0] coe_dat_wire242 = coe_dat_wire[2709:2700] ;
    wire [9:0] coe_dat_wire243 = coe_dat_wire[2699:2690] ;
    wire [9:0] coe_dat_wire244 = coe_dat_wire[2689:2680] ;
    wire [9:0] coe_dat_wire245 = coe_dat_wire[2679:2670] ;
    wire [9:0] coe_dat_wire246 = coe_dat_wire[2669:2660] ;
    wire [9:0] coe_dat_wire247 = coe_dat_wire[2659:2650] ;
    wire [9:0] coe_dat_wire248 = coe_dat_wire[2649:2640] ;
    wire [9:0] coe_dat_wire249 = coe_dat_wire[2639:2630] ;
    wire [9:0] coe_dat_wire250 = coe_dat_wire[2629:2620] ;
    wire [9:0] coe_dat_wire251 = coe_dat_wire[2619:2610] ;
    wire [9:0] coe_dat_wire252 = coe_dat_wire[2609:2600] ;
    wire [9:0] coe_dat_wire253 = coe_dat_wire[2599:2590] ;
    wire [9:0] coe_dat_wire254 = coe_dat_wire[2589:2580] ;
    wire [9:0] coe_dat_wire255 = coe_dat_wire[2579:2570] ;
    wire [9:0] coe_dat_wire256 = coe_dat_wire[2569:2560] ;
    wire [9:0] coe_dat_wire257 = coe_dat_wire[2559:2550] ;
    wire [9:0] coe_dat_wire258 = coe_dat_wire[2549:2540] ;
    wire [9:0] coe_dat_wire259 = coe_dat_wire[2539:2530] ;
    wire [9:0] coe_dat_wire260 = coe_dat_wire[2529:2520] ;
    wire [9:0] coe_dat_wire261 = coe_dat_wire[2519:2510] ;
    wire [9:0] coe_dat_wire262 = coe_dat_wire[2509:2500] ;
    wire [9:0] coe_dat_wire263 = coe_dat_wire[2499:2490] ;
    wire [9:0] coe_dat_wire264 = coe_dat_wire[2489:2480] ;
    wire [9:0] coe_dat_wire265 = coe_dat_wire[2479:2470] ;
    wire [9:0] coe_dat_wire266 = coe_dat_wire[2469:2460] ;
    wire [9:0] coe_dat_wire267 = coe_dat_wire[2459:2450] ;
    wire [9:0] coe_dat_wire268 = coe_dat_wire[2449:2440] ;
    wire [9:0] coe_dat_wire269 = coe_dat_wire[2439:2430] ;
    wire [9:0] coe_dat_wire270 = coe_dat_wire[2429:2420] ;
    wire [9:0] coe_dat_wire271 = coe_dat_wire[2419:2410] ;
    wire [9:0] coe_dat_wire272 = coe_dat_wire[2409:2400] ;
    wire [9:0] coe_dat_wire273 = coe_dat_wire[2399:2390] ;
    wire [9:0] coe_dat_wire274 = coe_dat_wire[2389:2380] ;
    wire [9:0] coe_dat_wire275 = coe_dat_wire[2379:2370] ;
    wire [9:0] coe_dat_wire276 = coe_dat_wire[2369:2360] ;
    wire [9:0] coe_dat_wire277 = coe_dat_wire[2359:2350] ;
    wire [9:0] coe_dat_wire278 = coe_dat_wire[2349:2340] ;
    wire [9:0] coe_dat_wire279 = coe_dat_wire[2339:2330] ;
    wire [9:0] coe_dat_wire280 = coe_dat_wire[2329:2320] ;
    wire [9:0] coe_dat_wire281 = coe_dat_wire[2319:2310] ;
    wire [9:0] coe_dat_wire282 = coe_dat_wire[2309:2300] ;
    wire [9:0] coe_dat_wire283 = coe_dat_wire[2299:2290] ;
    wire [9:0] coe_dat_wire284 = coe_dat_wire[2289:2280] ;
    wire [9:0] coe_dat_wire285 = coe_dat_wire[2279:2270] ;
    wire [9:0] coe_dat_wire286 = coe_dat_wire[2269:2260] ;
    wire [9:0] coe_dat_wire287 = coe_dat_wire[2259:2250] ;
    wire [9:0] coe_dat_wire288 = coe_dat_wire[2249:2240] ;
    wire [9:0] coe_dat_wire289 = coe_dat_wire[2239:2230] ;
    wire [9:0] coe_dat_wire290 = coe_dat_wire[2229:2220] ;
    wire [9:0] coe_dat_wire291 = coe_dat_wire[2219:2210] ;
    wire [9:0] coe_dat_wire292 = coe_dat_wire[2209:2200] ;
    wire [9:0] coe_dat_wire293 = coe_dat_wire[2199:2190] ;
    wire [9:0] coe_dat_wire294 = coe_dat_wire[2189:2180] ;
    wire [9:0] coe_dat_wire295 = coe_dat_wire[2179:2170] ;
    wire [9:0] coe_dat_wire296 = coe_dat_wire[2169:2160] ;
    wire [9:0] coe_dat_wire297 = coe_dat_wire[2159:2150] ;
    wire [9:0] coe_dat_wire298 = coe_dat_wire[2149:2140] ;
    wire [9:0] coe_dat_wire299 = coe_dat_wire[2139:2130] ;
    wire [9:0] coe_dat_wire300 = coe_dat_wire[2129:2120] ;
    wire [9:0] coe_dat_wire301 = coe_dat_wire[2119:2110] ;
    wire [9:0] coe_dat_wire302 = coe_dat_wire[2109:2100] ;
    wire [9:0] coe_dat_wire303 = coe_dat_wire[2099:2090] ;
    wire [9:0] coe_dat_wire304 = coe_dat_wire[2089:2080] ;
    wire [9:0] coe_dat_wire305 = coe_dat_wire[2079:2070] ;
    wire [9:0] coe_dat_wire306 = coe_dat_wire[2069:2060] ;
    wire [9:0] coe_dat_wire307 = coe_dat_wire[2059:2050] ;
    wire [9:0] coe_dat_wire308 = coe_dat_wire[2049:2040] ;
    wire [9:0] coe_dat_wire309 = coe_dat_wire[2039:2030] ;
    wire [9:0] coe_dat_wire310 = coe_dat_wire[2029:2020] ;
    wire [9:0] coe_dat_wire311 = coe_dat_wire[2019:2010] ;
    wire [9:0] coe_dat_wire312 = coe_dat_wire[2009:2000] ;
    wire [9:0] coe_dat_wire313 = coe_dat_wire[1999:1990] ;
    wire [9:0] coe_dat_wire314 = coe_dat_wire[1989:1980] ;
    wire [9:0] coe_dat_wire315 = coe_dat_wire[1979:1970] ;
    wire [9:0] coe_dat_wire316 = coe_dat_wire[1969:1960] ;
    wire [9:0] coe_dat_wire317 = coe_dat_wire[1959:1950] ;
    wire [9:0] coe_dat_wire318 = coe_dat_wire[1949:1940] ;
    wire [9:0] coe_dat_wire319 = coe_dat_wire[1939:1930] ;
    wire [9:0] coe_dat_wire320 = coe_dat_wire[1929:1920] ;
    wire [9:0] coe_dat_wire321 = coe_dat_wire[1919:1910] ;
    wire [9:0] coe_dat_wire322 = coe_dat_wire[1909:1900] ;
    wire [9:0] coe_dat_wire323 = coe_dat_wire[1899:1890] ;
    wire [9:0] coe_dat_wire324 = coe_dat_wire[1889:1880] ;
    wire [9:0] coe_dat_wire325 = coe_dat_wire[1879:1870] ;
    wire [9:0] coe_dat_wire326 = coe_dat_wire[1869:1860] ;
    wire [9:0] coe_dat_wire327 = coe_dat_wire[1859:1850] ;
    wire [9:0] coe_dat_wire328 = coe_dat_wire[1849:1840] ;
    wire [9:0] coe_dat_wire329 = coe_dat_wire[1839:1830] ;
    wire [9:0] coe_dat_wire330 = coe_dat_wire[1829:1820] ;
    wire [9:0] coe_dat_wire331 = coe_dat_wire[1819:1810] ;
    wire [9:0] coe_dat_wire332 = coe_dat_wire[1809:1800] ;
    wire [9:0] coe_dat_wire333 = coe_dat_wire[1799:1790] ;
    wire [9:0] coe_dat_wire334 = coe_dat_wire[1789:1780] ;
    wire [9:0] coe_dat_wire335 = coe_dat_wire[1779:1770] ;
    wire [9:0] coe_dat_wire336 = coe_dat_wire[1769:1760] ;
    wire [9:0] coe_dat_wire337 = coe_dat_wire[1759:1750] ;
    wire [9:0] coe_dat_wire338 = coe_dat_wire[1749:1740] ;
    wire [9:0] coe_dat_wire339 = coe_dat_wire[1739:1730] ;
    wire [9:0] coe_dat_wire340 = coe_dat_wire[1729:1720] ;
    wire [9:0] coe_dat_wire341 = coe_dat_wire[1719:1710] ;
    wire [9:0] coe_dat_wire342 = coe_dat_wire[1709:1700] ;
    wire [9:0] coe_dat_wire343 = coe_dat_wire[1699:1690] ;
    wire [9:0] coe_dat_wire344 = coe_dat_wire[1689:1680] ;
    wire [9:0] coe_dat_wire345 = coe_dat_wire[1679:1670] ;
    wire [9:0] coe_dat_wire346 = coe_dat_wire[1669:1660] ;
    wire [9:0] coe_dat_wire347 = coe_dat_wire[1659:1650] ;
    wire [9:0] coe_dat_wire348 = coe_dat_wire[1649:1640] ;
    wire [9:0] coe_dat_wire349 = coe_dat_wire[1639:1630] ;
    wire [9:0] coe_dat_wire350 = coe_dat_wire[1629:1620] ;
    wire [9:0] coe_dat_wire351 = coe_dat_wire[1619:1610] ;
    wire [9:0] coe_dat_wire352 = coe_dat_wire[1609:1600] ;
    wire [9:0] coe_dat_wire353 = coe_dat_wire[1599:1590] ;
    wire [9:0] coe_dat_wire354 = coe_dat_wire[1589:1580] ;
    wire [9:0] coe_dat_wire355 = coe_dat_wire[1579:1570] ;
    wire [9:0] coe_dat_wire356 = coe_dat_wire[1569:1560] ;
    wire [9:0] coe_dat_wire357 = coe_dat_wire[1559:1550] ;
    wire [9:0] coe_dat_wire358 = coe_dat_wire[1549:1540] ;
    wire [9:0] coe_dat_wire359 = coe_dat_wire[1539:1530] ;
    wire [9:0] coe_dat_wire360 = coe_dat_wire[1529:1520] ;
    wire [9:0] coe_dat_wire361 = coe_dat_wire[1519:1510] ;
    wire [9:0] coe_dat_wire362 = coe_dat_wire[1509:1500] ;
    wire [9:0] coe_dat_wire363 = coe_dat_wire[1499:1490] ;
    wire [9:0] coe_dat_wire364 = coe_dat_wire[1489:1480] ;
    wire [9:0] coe_dat_wire365 = coe_dat_wire[1479:1470] ;
    wire [9:0] coe_dat_wire366 = coe_dat_wire[1469:1460] ;
    wire [9:0] coe_dat_wire367 = coe_dat_wire[1459:1450] ;
    wire [9:0] coe_dat_wire368 = coe_dat_wire[1449:1440] ;
    wire [9:0] coe_dat_wire369 = coe_dat_wire[1439:1430] ;
    wire [9:0] coe_dat_wire370 = coe_dat_wire[1429:1420] ;
    wire [9:0] coe_dat_wire371 = coe_dat_wire[1419:1410] ;
    wire [9:0] coe_dat_wire372 = coe_dat_wire[1409:1400] ;
    wire [9:0] coe_dat_wire373 = coe_dat_wire[1399:1390] ;
    wire [9:0] coe_dat_wire374 = coe_dat_wire[1389:1380] ;
    wire [9:0] coe_dat_wire375 = coe_dat_wire[1379:1370] ;
    wire [9:0] coe_dat_wire376 = coe_dat_wire[1369:1360] ;
    wire [9:0] coe_dat_wire377 = coe_dat_wire[1359:1350] ;
    wire [9:0] coe_dat_wire378 = coe_dat_wire[1349:1340] ;
    wire [9:0] coe_dat_wire379 = coe_dat_wire[1339:1330] ;
    wire [9:0] coe_dat_wire380 = coe_dat_wire[1329:1320] ;
    wire [9:0] coe_dat_wire381 = coe_dat_wire[1319:1310] ;
    wire [9:0] coe_dat_wire382 = coe_dat_wire[1309:1300] ;
    wire [9:0] coe_dat_wire383 = coe_dat_wire[1299:1290] ;
    wire [9:0] coe_dat_wire384 = coe_dat_wire[1289:1280] ;
    wire [9:0] coe_dat_wire385 = coe_dat_wire[1279:1270] ;
    wire [9:0] coe_dat_wire386 = coe_dat_wire[1269:1260] ;
    wire [9:0] coe_dat_wire387 = coe_dat_wire[1259:1250] ;
    wire [9:0] coe_dat_wire388 = coe_dat_wire[1249:1240] ;
    wire [9:0] coe_dat_wire389 = coe_dat_wire[1239:1230] ;
    wire [9:0] coe_dat_wire390 = coe_dat_wire[1229:1220] ;
    wire [9:0] coe_dat_wire391 = coe_dat_wire[1219:1210] ;
    wire [9:0] coe_dat_wire392 = coe_dat_wire[1209:1200] ;
    wire [9:0] coe_dat_wire393 = coe_dat_wire[1199:1190] ;
    wire [9:0] coe_dat_wire394 = coe_dat_wire[1189:1180] ;
    wire [9:0] coe_dat_wire395 = coe_dat_wire[1179:1170] ;
    wire [9:0] coe_dat_wire396 = coe_dat_wire[1169:1160] ;
    wire [9:0] coe_dat_wire397 = coe_dat_wire[1159:1150] ;
    wire [9:0] coe_dat_wire398 = coe_dat_wire[1149:1140] ;
    wire [9:0] coe_dat_wire399 = coe_dat_wire[1139:1130] ;
    wire [9:0] coe_dat_wire400 = coe_dat_wire[1129:1120] ;
    wire [9:0] coe_dat_wire401 = coe_dat_wire[1119:1110] ;
    wire [9:0] coe_dat_wire402 = coe_dat_wire[1109:1100] ;
    wire [9:0] coe_dat_wire403 = coe_dat_wire[1099:1090] ;
    wire [9:0] coe_dat_wire404 = coe_dat_wire[1089:1080] ;
    wire [9:0] coe_dat_wire405 = coe_dat_wire[1079:1070] ;
    wire [9:0] coe_dat_wire406 = coe_dat_wire[1069:1060] ;
    wire [9:0] coe_dat_wire407 = coe_dat_wire[1059:1050] ;
    wire [9:0] coe_dat_wire408 = coe_dat_wire[1049:1040] ;
    wire [9:0] coe_dat_wire409 = coe_dat_wire[1039:1030] ;
    wire [9:0] coe_dat_wire410 = coe_dat_wire[1029:1020] ;
    wire [9:0] coe_dat_wire411 = coe_dat_wire[1019:1010] ;
    wire [9:0] coe_dat_wire412 = coe_dat_wire[1009:1000] ;
    wire [9:0] coe_dat_wire413 = coe_dat_wire[999:990] ;
    wire [9:0] coe_dat_wire414 = coe_dat_wire[989:980] ;
    wire [9:0] coe_dat_wire415 = coe_dat_wire[979:970] ;
    wire [9:0] coe_dat_wire416 = coe_dat_wire[969:960] ;
    wire [9:0] coe_dat_wire417 = coe_dat_wire[959:950] ;
    wire [9:0] coe_dat_wire418 = coe_dat_wire[949:940] ;
    wire [9:0] coe_dat_wire419 = coe_dat_wire[939:930] ;
    wire [9:0] coe_dat_wire420 = coe_dat_wire[929:920] ;
    wire [9:0] coe_dat_wire421 = coe_dat_wire[919:910] ;
    wire [9:0] coe_dat_wire422 = coe_dat_wire[909:900] ;
    wire [9:0] coe_dat_wire423 = coe_dat_wire[899:890] ;
    wire [9:0] coe_dat_wire424 = coe_dat_wire[889:880] ;
    wire [9:0] coe_dat_wire425 = coe_dat_wire[879:870] ;
    wire [9:0] coe_dat_wire426 = coe_dat_wire[869:860] ;
    wire [9:0] coe_dat_wire427 = coe_dat_wire[859:850] ;
    wire [9:0] coe_dat_wire428 = coe_dat_wire[849:840] ;
    wire [9:0] coe_dat_wire429 = coe_dat_wire[839:830] ;
    wire [9:0] coe_dat_wire430 = coe_dat_wire[829:820] ;
    wire [9:0] coe_dat_wire431 = coe_dat_wire[819:810] ;
    wire [9:0] coe_dat_wire432 = coe_dat_wire[809:800] ;
    wire [9:0] coe_dat_wire433 = coe_dat_wire[799:790] ;
    wire [9:0] coe_dat_wire434 = coe_dat_wire[789:780] ;
    wire [9:0] coe_dat_wire435 = coe_dat_wire[779:770] ;
    wire [9:0] coe_dat_wire436 = coe_dat_wire[769:760] ;
    wire [9:0] coe_dat_wire437 = coe_dat_wire[759:750] ;
    wire [9:0] coe_dat_wire438 = coe_dat_wire[749:740] ;
    wire [9:0] coe_dat_wire439 = coe_dat_wire[739:730] ;
    wire [9:0] coe_dat_wire440 = coe_dat_wire[729:720] ;
    wire [9:0] coe_dat_wire441 = coe_dat_wire[719:710] ;
    wire [9:0] coe_dat_wire442 = coe_dat_wire[709:700] ;
    wire [9:0] coe_dat_wire443 = coe_dat_wire[699:690] ;
    wire [9:0] coe_dat_wire444 = coe_dat_wire[689:680] ;
    wire [9:0] coe_dat_wire445 = coe_dat_wire[679:670] ;
    wire [9:0] coe_dat_wire446 = coe_dat_wire[669:660] ;
    wire [9:0] coe_dat_wire447 = coe_dat_wire[659:650] ;
    wire [9:0] coe_dat_wire448 = coe_dat_wire[649:640] ;
    wire [9:0] coe_dat_wire449 = coe_dat_wire[639:630] ;
    wire [9:0] coe_dat_wire450 = coe_dat_wire[629:620] ;
    wire [9:0] coe_dat_wire451 = coe_dat_wire[619:610] ;
    wire [9:0] coe_dat_wire452 = coe_dat_wire[609:600] ;
    wire [9:0] coe_dat_wire453 = coe_dat_wire[599:590] ;
    wire [9:0] coe_dat_wire454 = coe_dat_wire[589:580] ;
    wire [9:0] coe_dat_wire455 = coe_dat_wire[579:570] ;
    wire [9:0] coe_dat_wire456 = coe_dat_wire[569:560] ;
    wire [9:0] coe_dat_wire457 = coe_dat_wire[559:550] ;
    wire [9:0] coe_dat_wire458 = coe_dat_wire[549:540] ;
    wire [9:0] coe_dat_wire459 = coe_dat_wire[539:530] ;
    wire [9:0] coe_dat_wire460 = coe_dat_wire[529:520] ;
    wire [9:0] coe_dat_wire461 = coe_dat_wire[519:510] ;
    wire [9:0] coe_dat_wire462 = coe_dat_wire[509:500] ;
    wire [9:0] coe_dat_wire463 = coe_dat_wire[499:490] ;
    wire [9:0] coe_dat_wire464 = coe_dat_wire[489:480] ;
    wire [9:0] coe_dat_wire465 = coe_dat_wire[479:470] ;
    wire [9:0] coe_dat_wire466 = coe_dat_wire[469:460] ;
    wire [9:0] coe_dat_wire467 = coe_dat_wire[459:450] ;
    wire [9:0] coe_dat_wire468 = coe_dat_wire[449:440] ;
    wire [9:0] coe_dat_wire469 = coe_dat_wire[439:430] ;
    wire [9:0] coe_dat_wire470 = coe_dat_wire[429:420] ;
    wire [9:0] coe_dat_wire471 = coe_dat_wire[419:410] ;
    wire [9:0] coe_dat_wire472 = coe_dat_wire[409:400] ;
    wire [9:0] coe_dat_wire473 = coe_dat_wire[399:390] ;
    wire [9:0] coe_dat_wire474 = coe_dat_wire[389:380] ;
    wire [9:0] coe_dat_wire475 = coe_dat_wire[379:370] ;
    wire [9:0] coe_dat_wire476 = coe_dat_wire[369:360] ;
    wire [9:0] coe_dat_wire477 = coe_dat_wire[359:350] ;
    wire [9:0] coe_dat_wire478 = coe_dat_wire[349:340] ;
    wire [9:0] coe_dat_wire479 = coe_dat_wire[339:330] ;
    wire [9:0] coe_dat_wire480 = coe_dat_wire[329:320] ;
    wire [9:0] coe_dat_wire481 = coe_dat_wire[319:310] ;
    wire [9:0] coe_dat_wire482 = coe_dat_wire[309:300] ;
    wire [9:0] coe_dat_wire483 = coe_dat_wire[299:290] ;
    wire [9:0] coe_dat_wire484 = coe_dat_wire[289:280] ;
    wire [9:0] coe_dat_wire485 = coe_dat_wire[279:270] ;
    wire [9:0] coe_dat_wire486 = coe_dat_wire[269:260] ;
    wire [9:0] coe_dat_wire487 = coe_dat_wire[259:250] ;
    wire [9:0] coe_dat_wire488 = coe_dat_wire[249:240] ;
    wire [9:0] coe_dat_wire489 = coe_dat_wire[239:230] ;
    wire [9:0] coe_dat_wire490 = coe_dat_wire[229:220] ;
    wire [9:0] coe_dat_wire491 = coe_dat_wire[219:210] ;
    wire [9:0] coe_dat_wire492 = coe_dat_wire[209:200] ;
    wire [9:0] coe_dat_wire493 = coe_dat_wire[199:190] ;
    wire [9:0] coe_dat_wire494 = coe_dat_wire[189:180] ;
    wire [9:0] coe_dat_wire495 = coe_dat_wire[179:170] ;
    wire [9:0] coe_dat_wire496 = coe_dat_wire[169:160] ;
    wire [9:0] coe_dat_wire497 = coe_dat_wire[159:150] ;
    wire [9:0] coe_dat_wire498 = coe_dat_wire[149:140] ;
    wire [9:0] coe_dat_wire499 = coe_dat_wire[139:130] ;
    wire [9:0] coe_dat_wire500 = coe_dat_wire[129:120] ;
    wire [9:0] coe_dat_wire501 = coe_dat_wire[119:110] ;
    wire [9:0] coe_dat_wire502 = coe_dat_wire[109:100] ;
    wire [9:0] coe_dat_wire503 = coe_dat_wire[99:90] ;
    wire [9:0] coe_dat_wire504 = coe_dat_wire[89:80] ;
    wire [9:0] coe_dat_wire505 = coe_dat_wire[79:70] ;
    wire [9:0] coe_dat_wire506 = coe_dat_wire[69:60] ;
    wire [9:0] coe_dat_wire507 = coe_dat_wire[59:50] ;
    wire [9:0] coe_dat_wire508 = coe_dat_wire[49:40] ;
    wire [9:0] coe_dat_wire509 = coe_dat_wire[39:30] ;
    wire [9:0] coe_dat_wire510 = coe_dat_wire[29:20] ;
    wire [9:0] coe_dat_wire511 = coe_dat_wire[19:10] ;
    wire [9:0] coe_dat_wire512 = coe_dat_wire[9:0] ;
                                                 
    reg [9:0] in_dat_hld01,  in_dat_hld02,  in_dat_hld03,  in_dat_hld04,  in_dat_hld05,  in_dat_hld06,  in_dat_hld07,  in_dat_hld08,
              in_dat_hld09,  in_dat_hld10,  in_dat_hld11,  in_dat_hld12,  in_dat_hld13,  in_dat_hld14,  in_dat_hld15,  in_dat_hld16,
              in_dat_hld17,  in_dat_hld18,  in_dat_hld19,  in_dat_hld20,  in_dat_hld21,  in_dat_hld22,  in_dat_hld23,  in_dat_hld24,
              in_dat_hld25,  in_dat_hld26,  in_dat_hld27,  in_dat_hld28,  in_dat_hld29,  in_dat_hld30,  in_dat_hld31,  in_dat_hld32,
              in_dat_hld33,  in_dat_hld34,  in_dat_hld35,  in_dat_hld36,  in_dat_hld37,  in_dat_hld38,  in_dat_hld39,  in_dat_hld40,
              in_dat_hld41,  in_dat_hld42,  in_dat_hld43,  in_dat_hld44,  in_dat_hld45,  in_dat_hld46,  in_dat_hld47,  in_dat_hld48,
              in_dat_hld49,  in_dat_hld50,  in_dat_hld51,  in_dat_hld52,  in_dat_hld53,  in_dat_hld54,  in_dat_hld55,  in_dat_hld56,
              in_dat_hld57,  in_dat_hld58,  in_dat_hld59,  in_dat_hld60,  in_dat_hld61,  in_dat_hld62,  in_dat_hld63,  in_dat_hld64,
              in_dat_hld65,  in_dat_hld66,  in_dat_hld67,  in_dat_hld68,  in_dat_hld69,  in_dat_hld70,  in_dat_hld71,  in_dat_hld72,
              in_dat_hld73,  in_dat_hld74,  in_dat_hld75,  in_dat_hld76,  in_dat_hld77,  in_dat_hld78,  in_dat_hld79,  in_dat_hld80,
              in_dat_hld81,  in_dat_hld82,  in_dat_hld83,  in_dat_hld84,  in_dat_hld85,  in_dat_hld86,  in_dat_hld87,  in_dat_hld88,
              in_dat_hld89,  in_dat_hld90,  in_dat_hld91,  in_dat_hld92,  in_dat_hld93,  in_dat_hld94,  in_dat_hld95,  in_dat_hld96,
              in_dat_hld97,  in_dat_hld98,  in_dat_hld99,  in_dat_hld100, in_dat_hld101, in_dat_hld102, in_dat_hld103, in_dat_hld104,
              in_dat_hld105, in_dat_hld106, in_dat_hld107, in_dat_hld108, in_dat_hld109, in_dat_hld110, in_dat_hld111, in_dat_hld112,
              in_dat_hld113, in_dat_hld114, in_dat_hld115, in_dat_hld116, in_dat_hld117, in_dat_hld118, in_dat_hld119, in_dat_hld120,
              in_dat_hld121, in_dat_hld122, in_dat_hld123, in_dat_hld124, in_dat_hld125, in_dat_hld126, in_dat_hld127, in_dat_hld128,
              in_dat_hld129, in_dat_hld130, in_dat_hld131, in_dat_hld132, in_dat_hld133, in_dat_hld134, in_dat_hld135, in_dat_hld136,
              in_dat_hld137, in_dat_hld138, in_dat_hld139, in_dat_hld140, in_dat_hld141, in_dat_hld142, in_dat_hld143, in_dat_hld144,
              in_dat_hld145, in_dat_hld146, in_dat_hld147, in_dat_hld148, in_dat_hld149, in_dat_hld150, in_dat_hld151, in_dat_hld152,
              in_dat_hld153, in_dat_hld154, in_dat_hld155, in_dat_hld156, in_dat_hld157, in_dat_hld158, in_dat_hld159, in_dat_hld160,
              in_dat_hld161, in_dat_hld162, in_dat_hld163, in_dat_hld164, in_dat_hld165, in_dat_hld166, in_dat_hld167, in_dat_hld168,
              in_dat_hld169, in_dat_hld170, in_dat_hld171, in_dat_hld172, in_dat_hld173, in_dat_hld174, in_dat_hld175, in_dat_hld176,
              in_dat_hld177, in_dat_hld178, in_dat_hld179, in_dat_hld180, in_dat_hld181, in_dat_hld182, in_dat_hld183, in_dat_hld184,
              in_dat_hld185, in_dat_hld186, in_dat_hld187, in_dat_hld188, in_dat_hld189, in_dat_hld190, in_dat_hld191, in_dat_hld192,
              in_dat_hld193, in_dat_hld194, in_dat_hld195, in_dat_hld196, in_dat_hld197, in_dat_hld198, in_dat_hld199, in_dat_hld200,
              in_dat_hld201, in_dat_hld202, in_dat_hld203, in_dat_hld204, in_dat_hld205, in_dat_hld206, in_dat_hld207, in_dat_hld208,
              in_dat_hld209, in_dat_hld210, in_dat_hld211, in_dat_hld212, in_dat_hld213, in_dat_hld214, in_dat_hld215, in_dat_hld216,
              in_dat_hld217, in_dat_hld218, in_dat_hld219, in_dat_hld220, in_dat_hld221, in_dat_hld222, in_dat_hld223, in_dat_hld224,
              in_dat_hld225, in_dat_hld226, in_dat_hld227, in_dat_hld228, in_dat_hld229, in_dat_hld230, in_dat_hld231, in_dat_hld232,
              in_dat_hld233, in_dat_hld234, in_dat_hld235, in_dat_hld236, in_dat_hld237, in_dat_hld238, in_dat_hld239, in_dat_hld240,
              in_dat_hld241, in_dat_hld242, in_dat_hld243, in_dat_hld244, in_dat_hld245, in_dat_hld246, in_dat_hld247, in_dat_hld248,
              in_dat_hld249, in_dat_hld250, in_dat_hld251, in_dat_hld252, in_dat_hld253, in_dat_hld254, in_dat_hld255, in_dat_hld256,
              in_dat_hld257, in_dat_hld258, in_dat_hld259, in_dat_hld260, in_dat_hld261, in_dat_hld262, in_dat_hld263, in_dat_hld264,
              in_dat_hld265, in_dat_hld266, in_dat_hld267, in_dat_hld268, in_dat_hld269, in_dat_hld270, in_dat_hld271, in_dat_hld272,
              in_dat_hld273, in_dat_hld274, in_dat_hld275, in_dat_hld276, in_dat_hld277, in_dat_hld278, in_dat_hld279, in_dat_hld280,
              in_dat_hld281, in_dat_hld282, in_dat_hld283, in_dat_hld284, in_dat_hld285, in_dat_hld286, in_dat_hld287, in_dat_hld288,
              in_dat_hld289, in_dat_hld290, in_dat_hld291, in_dat_hld292, in_dat_hld293, in_dat_hld294, in_dat_hld295, in_dat_hld296,
              in_dat_hld297, in_dat_hld298, in_dat_hld299, in_dat_hld300, in_dat_hld301, in_dat_hld302, in_dat_hld303, in_dat_hld304,
              in_dat_hld305, in_dat_hld306, in_dat_hld307, in_dat_hld308, in_dat_hld309, in_dat_hld310, in_dat_hld311, in_dat_hld312,
              in_dat_hld313, in_dat_hld314, in_dat_hld315, in_dat_hld316, in_dat_hld317, in_dat_hld318, in_dat_hld319, in_dat_hld320,
              in_dat_hld321, in_dat_hld322, in_dat_hld323, in_dat_hld324, in_dat_hld325, in_dat_hld326, in_dat_hld327, in_dat_hld328,
              in_dat_hld329, in_dat_hld330, in_dat_hld331, in_dat_hld332, in_dat_hld333, in_dat_hld334, in_dat_hld335, in_dat_hld336,
              in_dat_hld337, in_dat_hld338, in_dat_hld339, in_dat_hld340, in_dat_hld341, in_dat_hld342, in_dat_hld343, in_dat_hld344,
              in_dat_hld345, in_dat_hld346, in_dat_hld347, in_dat_hld348, in_dat_hld349, in_dat_hld350, in_dat_hld351, in_dat_hld352,
              in_dat_hld353, in_dat_hld354, in_dat_hld355, in_dat_hld356, in_dat_hld357, in_dat_hld358, in_dat_hld359, in_dat_hld360,
              in_dat_hld361, in_dat_hld362, in_dat_hld363, in_dat_hld364, in_dat_hld365, in_dat_hld366, in_dat_hld367, in_dat_hld368,
              in_dat_hld369, in_dat_hld370, in_dat_hld371, in_dat_hld372, in_dat_hld373, in_dat_hld374, in_dat_hld375, in_dat_hld376,
              in_dat_hld377, in_dat_hld378, in_dat_hld379, in_dat_hld380, in_dat_hld381, in_dat_hld382, in_dat_hld383, in_dat_hld384,
              in_dat_hld385, in_dat_hld386, in_dat_hld387, in_dat_hld388, in_dat_hld389, in_dat_hld390, in_dat_hld391, in_dat_hld392,
              in_dat_hld393, in_dat_hld394, in_dat_hld395, in_dat_hld396, in_dat_hld397, in_dat_hld398, in_dat_hld399, in_dat_hld400,
              in_dat_hld401, in_dat_hld402, in_dat_hld403, in_dat_hld404, in_dat_hld405, in_dat_hld406, in_dat_hld407, in_dat_hld408,
              in_dat_hld409, in_dat_hld410, in_dat_hld411, in_dat_hld412, in_dat_hld413, in_dat_hld414, in_dat_hld415, in_dat_hld416,
              in_dat_hld417, in_dat_hld418, in_dat_hld419, in_dat_hld420, in_dat_hld421, in_dat_hld422, in_dat_hld423, in_dat_hld424,
              in_dat_hld425, in_dat_hld426, in_dat_hld427, in_dat_hld428, in_dat_hld429, in_dat_hld430, in_dat_hld431, in_dat_hld432,
              in_dat_hld433, in_dat_hld434, in_dat_hld435, in_dat_hld436, in_dat_hld437, in_dat_hld438, in_dat_hld439, in_dat_hld440,
              in_dat_hld441, in_dat_hld442, in_dat_hld443, in_dat_hld444, in_dat_hld445, in_dat_hld446, in_dat_hld447, in_dat_hld448,
              in_dat_hld449, in_dat_hld450, in_dat_hld451, in_dat_hld452, in_dat_hld453, in_dat_hld454, in_dat_hld455, in_dat_hld456,
              in_dat_hld457, in_dat_hld458, in_dat_hld459, in_dat_hld460, in_dat_hld461, in_dat_hld462, in_dat_hld463, in_dat_hld464,
              in_dat_hld465, in_dat_hld466, in_dat_hld467, in_dat_hld468, in_dat_hld469, in_dat_hld470, in_dat_hld471, in_dat_hld472,
              in_dat_hld473, in_dat_hld474, in_dat_hld475, in_dat_hld476, in_dat_hld477, in_dat_hld478, in_dat_hld479, in_dat_hld480,
              in_dat_hld481, in_dat_hld482, in_dat_hld483, in_dat_hld484, in_dat_hld485, in_dat_hld486, in_dat_hld487, in_dat_hld488,
              in_dat_hld489, in_dat_hld490, in_dat_hld491, in_dat_hld492, in_dat_hld493, in_dat_hld494, in_dat_hld495, in_dat_hld496,
              in_dat_hld497, in_dat_hld498, in_dat_hld499, in_dat_hld500, in_dat_hld501, in_dat_hld502, in_dat_hld503, in_dat_hld504,
              in_dat_hld505, in_dat_hld506, in_dat_hld507, in_dat_hld508, in_dat_hld509, in_dat_hld510, in_dat_hld511, in_dat_hld512; 

    always @ (posedge clk) begin
		if(rst) begin
            in_dat_hld01[9:0]  <= #DLY 10'd0 ;
            in_dat_hld02[9:0]  <= #DLY 10'd0 ;
            in_dat_hld03[9:0]  <= #DLY 10'd0 ;
            in_dat_hld04[9:0]  <= #DLY 10'd0 ;
            in_dat_hld05[9:0]  <= #DLY 10'd0 ;
            in_dat_hld06[9:0]  <= #DLY 10'd0 ;
            in_dat_hld07[9:0]  <= #DLY 10'd0 ;
            in_dat_hld08[9:0]  <= #DLY 10'd0 ;
            in_dat_hld09[9:0]  <= #DLY 10'd0 ;
            in_dat_hld10[9:0]  <= #DLY 10'd0 ;
            in_dat_hld11[9:0]  <= #DLY 10'd0 ;
            in_dat_hld12[9:0]  <= #DLY 10'd0 ;
            in_dat_hld13[9:0]  <= #DLY 10'd0 ;
            in_dat_hld14[9:0]  <= #DLY 10'd0 ;
            in_dat_hld15[9:0]  <= #DLY 10'd0 ;
            in_dat_hld16[9:0]  <= #DLY 10'd0 ;
            in_dat_hld17[9:0]  <= #DLY 10'd0 ;
            in_dat_hld18[9:0]  <= #DLY 10'd0 ;
            in_dat_hld19[9:0]  <= #DLY 10'd0 ;
            in_dat_hld20[9:0]  <= #DLY 10'd0 ;
            in_dat_hld21[9:0]  <= #DLY 10'd0 ;
            in_dat_hld22[9:0]  <= #DLY 10'd0 ;
            in_dat_hld23[9:0]  <= #DLY 10'd0 ;
            in_dat_hld24[9:0]  <= #DLY 10'd0 ;
            in_dat_hld25[9:0]  <= #DLY 10'd0 ;
            in_dat_hld26[9:0]  <= #DLY 10'd0 ;
            in_dat_hld27[9:0]  <= #DLY 10'd0 ;
            in_dat_hld28[9:0]  <= #DLY 10'd0 ;
            in_dat_hld29[9:0]  <= #DLY 10'd0 ;
            in_dat_hld30[9:0]  <= #DLY 10'd0 ;
            in_dat_hld31[9:0]  <= #DLY 10'd0 ;
            in_dat_hld32[9:0]  <= #DLY 10'd0 ;
            in_dat_hld33[9:0]  <= #DLY 10'd0 ;
            in_dat_hld34[9:0]  <= #DLY 10'd0 ;
            in_dat_hld35[9:0]  <= #DLY 10'd0 ;
            in_dat_hld36[9:0]  <= #DLY 10'd0 ;
            in_dat_hld37[9:0]  <= #DLY 10'd0 ;
            in_dat_hld38[9:0]  <= #DLY 10'd0 ;
            in_dat_hld39[9:0]  <= #DLY 10'd0 ;
            in_dat_hld40[9:0]  <= #DLY 10'd0 ;
            in_dat_hld41[9:0]  <= #DLY 10'd0 ;
            in_dat_hld42[9:0]  <= #DLY 10'd0 ;
            in_dat_hld43[9:0]  <= #DLY 10'd0 ;
            in_dat_hld44[9:0]  <= #DLY 10'd0 ;
            in_dat_hld45[9:0]  <= #DLY 10'd0 ;
            in_dat_hld46[9:0]  <= #DLY 10'd0 ;
            in_dat_hld47[9:0]  <= #DLY 10'd0 ;
            in_dat_hld48[9:0]  <= #DLY 10'd0 ;
            in_dat_hld49[9:0]  <= #DLY 10'd0 ;
            in_dat_hld50[9:0]  <= #DLY 10'd0 ;
            in_dat_hld51[9:0]  <= #DLY 10'd0 ;
            in_dat_hld52[9:0]  <= #DLY 10'd0 ;
            in_dat_hld53[9:0]  <= #DLY 10'd0 ;
            in_dat_hld54[9:0]  <= #DLY 10'd0 ;
            in_dat_hld55[9:0]  <= #DLY 10'd0 ;
            in_dat_hld56[9:0]  <= #DLY 10'd0 ;
            in_dat_hld57[9:0]  <= #DLY 10'd0 ;
            in_dat_hld58[9:0]  <= #DLY 10'd0 ;
            in_dat_hld59[9:0]  <= #DLY 10'd0 ;
            in_dat_hld60[9:0]  <= #DLY 10'd0 ;
            in_dat_hld61[9:0]  <= #DLY 10'd0 ;
            in_dat_hld62[9:0]  <= #DLY 10'd0 ;
            in_dat_hld63[9:0]  <= #DLY 10'd0 ;
            in_dat_hld64[9:0]  <= #DLY 10'd0 ;
            in_dat_hld65[9:0]  <= #DLY 10'd0 ;
            in_dat_hld66[9:0]  <= #DLY 10'd0 ;
            in_dat_hld67[9:0]  <= #DLY 10'd0 ;
            in_dat_hld68[9:0]  <= #DLY 10'd0 ;
            in_dat_hld69[9:0]  <= #DLY 10'd0 ;
            in_dat_hld70[9:0]  <= #DLY 10'd0 ;
            in_dat_hld71[9:0]  <= #DLY 10'd0 ;
            in_dat_hld72[9:0]  <= #DLY 10'd0 ;
            in_dat_hld73[9:0]  <= #DLY 10'd0 ;
            in_dat_hld74[9:0]  <= #DLY 10'd0 ;
            in_dat_hld75[9:0]  <= #DLY 10'd0 ;
            in_dat_hld76[9:0]  <= #DLY 10'd0 ;
            in_dat_hld77[9:0]  <= #DLY 10'd0 ;
            in_dat_hld78[9:0]  <= #DLY 10'd0 ;
            in_dat_hld79[9:0]  <= #DLY 10'd0 ;
            in_dat_hld80[9:0]  <= #DLY 10'd0 ;
            in_dat_hld81[9:0]  <= #DLY 10'd0 ;
            in_dat_hld82[9:0]  <= #DLY 10'd0 ;
            in_dat_hld83[9:0]  <= #DLY 10'd0 ;
            in_dat_hld84[9:0]  <= #DLY 10'd0 ;
            in_dat_hld85[9:0]  <= #DLY 10'd0 ;
            in_dat_hld86[9:0]  <= #DLY 10'd0 ;
            in_dat_hld87[9:0]  <= #DLY 10'd0 ;
            in_dat_hld88[9:0]  <= #DLY 10'd0 ;
            in_dat_hld89[9:0]  <= #DLY 10'd0 ;
            in_dat_hld90[9:0]  <= #DLY 10'd0 ;
            in_dat_hld91[9:0]  <= #DLY 10'd0 ;
            in_dat_hld92[9:0]  <= #DLY 10'd0 ;
            in_dat_hld93[9:0]  <= #DLY 10'd0 ;
            in_dat_hld94[9:0]  <= #DLY 10'd0 ;
            in_dat_hld95[9:0]  <= #DLY 10'd0 ;
            in_dat_hld96[9:0]  <= #DLY 10'd0 ;
            in_dat_hld97[9:0]  <= #DLY 10'd0 ;
            in_dat_hld98[9:0]  <= #DLY 10'd0 ;
            in_dat_hld99[9:0]  <= #DLY 10'd0 ;
            in_dat_hld100[9:0] <= #DLY 10'd0 ;
            in_dat_hld101[9:0] <= #DLY 10'd0 ;
            in_dat_hld102[9:0] <= #DLY 10'd0 ;
            in_dat_hld103[9:0] <= #DLY 10'd0 ;
            in_dat_hld104[9:0] <= #DLY 10'd0 ;
            in_dat_hld105[9:0] <= #DLY 10'd0 ;
            in_dat_hld106[9:0] <= #DLY 10'd0 ;
            in_dat_hld107[9:0] <= #DLY 10'd0 ;
            in_dat_hld108[9:0] <= #DLY 10'd0 ;
            in_dat_hld109[9:0] <= #DLY 10'd0 ;
            in_dat_hld110[9:0] <= #DLY 10'd0 ;
            in_dat_hld111[9:0] <= #DLY 10'd0 ;
            in_dat_hld112[9:0] <= #DLY 10'd0 ;
            in_dat_hld113[9:0] <= #DLY 10'd0 ;
            in_dat_hld114[9:0] <= #DLY 10'd0 ;
            in_dat_hld115[9:0] <= #DLY 10'd0 ;
            in_dat_hld116[9:0] <= #DLY 10'd0 ;
            in_dat_hld117[9:0] <= #DLY 10'd0 ;
            in_dat_hld118[9:0] <= #DLY 10'd0 ;
            in_dat_hld119[9:0] <= #DLY 10'd0 ;
            in_dat_hld120[9:0] <= #DLY 10'd0 ;
            in_dat_hld121[9:0] <= #DLY 10'd0 ;
            in_dat_hld122[9:0] <= #DLY 10'd0 ;
            in_dat_hld123[9:0] <= #DLY 10'd0 ;
            in_dat_hld124[9:0] <= #DLY 10'd0 ;
            in_dat_hld125[9:0] <= #DLY 10'd0 ;
            in_dat_hld126[9:0] <= #DLY 10'd0 ;
            in_dat_hld127[9:0] <= #DLY 10'd0 ;
            in_dat_hld128[9:0] <= #DLY 10'd0 ;
            in_dat_hld129[9:0] <= #DLY 10'd0 ;
            in_dat_hld130[9:0] <= #DLY 10'd0 ;
            in_dat_hld131[9:0] <= #DLY 10'd0 ;
            in_dat_hld132[9:0] <= #DLY 10'd0 ;
            in_dat_hld133[9:0] <= #DLY 10'd0 ;
            in_dat_hld134[9:0] <= #DLY 10'd0 ;
            in_dat_hld135[9:0] <= #DLY 10'd0 ;
            in_dat_hld136[9:0] <= #DLY 10'd0 ;
            in_dat_hld137[9:0] <= #DLY 10'd0 ;
            in_dat_hld138[9:0] <= #DLY 10'd0 ;
            in_dat_hld139[9:0] <= #DLY 10'd0 ;
            in_dat_hld140[9:0] <= #DLY 10'd0 ;
            in_dat_hld141[9:0] <= #DLY 10'd0 ;
            in_dat_hld142[9:0] <= #DLY 10'd0 ;
            in_dat_hld143[9:0] <= #DLY 10'd0 ;
            in_dat_hld144[9:0] <= #DLY 10'd0 ;
            in_dat_hld145[9:0] <= #DLY 10'd0 ;
            in_dat_hld146[9:0] <= #DLY 10'd0 ;
            in_dat_hld147[9:0] <= #DLY 10'd0 ;
            in_dat_hld148[9:0] <= #DLY 10'd0 ;
            in_dat_hld149[9:0] <= #DLY 10'd0 ;
            in_dat_hld150[9:0] <= #DLY 10'd0 ;
            in_dat_hld151[9:0] <= #DLY 10'd0 ;
            in_dat_hld152[9:0] <= #DLY 10'd0 ;
            in_dat_hld153[9:0] <= #DLY 10'd0 ;
            in_dat_hld154[9:0] <= #DLY 10'd0 ;
            in_dat_hld155[9:0] <= #DLY 10'd0 ;
            in_dat_hld156[9:0] <= #DLY 10'd0 ;
            in_dat_hld157[9:0] <= #DLY 10'd0 ;
            in_dat_hld158[9:0] <= #DLY 10'd0 ;
            in_dat_hld159[9:0] <= #DLY 10'd0 ;
            in_dat_hld160[9:0] <= #DLY 10'd0 ;
            in_dat_hld161[9:0] <= #DLY 10'd0 ;
            in_dat_hld162[9:0] <= #DLY 10'd0 ;
            in_dat_hld163[9:0] <= #DLY 10'd0 ;
            in_dat_hld164[9:0] <= #DLY 10'd0 ;
            in_dat_hld165[9:0] <= #DLY 10'd0 ;
            in_dat_hld166[9:0] <= #DLY 10'd0 ;
            in_dat_hld167[9:0] <= #DLY 10'd0 ;
            in_dat_hld168[9:0] <= #DLY 10'd0 ;
            in_dat_hld169[9:0] <= #DLY 10'd0 ;
            in_dat_hld170[9:0] <= #DLY 10'd0 ;
            in_dat_hld171[9:0] <= #DLY 10'd0 ;
            in_dat_hld172[9:0] <= #DLY 10'd0 ;
            in_dat_hld173[9:0] <= #DLY 10'd0 ;
            in_dat_hld174[9:0] <= #DLY 10'd0 ;
            in_dat_hld175[9:0] <= #DLY 10'd0 ;
            in_dat_hld176[9:0] <= #DLY 10'd0 ;
            in_dat_hld177[9:0] <= #DLY 10'd0 ;
            in_dat_hld178[9:0] <= #DLY 10'd0 ;
            in_dat_hld179[9:0] <= #DLY 10'd0 ;
            in_dat_hld180[9:0] <= #DLY 10'd0 ;
            in_dat_hld181[9:0] <= #DLY 10'd0 ;
            in_dat_hld182[9:0] <= #DLY 10'd0 ;
            in_dat_hld183[9:0] <= #DLY 10'd0 ;
            in_dat_hld184[9:0] <= #DLY 10'd0 ;
            in_dat_hld185[9:0] <= #DLY 10'd0 ;
            in_dat_hld186[9:0] <= #DLY 10'd0 ;
            in_dat_hld187[9:0] <= #DLY 10'd0 ;
            in_dat_hld188[9:0] <= #DLY 10'd0 ;
            in_dat_hld189[9:0] <= #DLY 10'd0 ;
            in_dat_hld190[9:0] <= #DLY 10'd0 ;
            in_dat_hld191[9:0] <= #DLY 10'd0 ;
            in_dat_hld192[9:0] <= #DLY 10'd0 ;
            in_dat_hld193[9:0] <= #DLY 10'd0 ;
            in_dat_hld194[9:0] <= #DLY 10'd0 ;
            in_dat_hld195[9:0] <= #DLY 10'd0 ;
            in_dat_hld196[9:0] <= #DLY 10'd0 ;
            in_dat_hld197[9:0] <= #DLY 10'd0 ;
            in_dat_hld198[9:0] <= #DLY 10'd0 ;
            in_dat_hld199[9:0] <= #DLY 10'd0 ;
            in_dat_hld200[9:0] <= #DLY 10'd0 ;
            in_dat_hld201[9:0] <= #DLY 10'd0 ;
            in_dat_hld202[9:0] <= #DLY 10'd0 ;
            in_dat_hld203[9:0] <= #DLY 10'd0 ;
            in_dat_hld204[9:0] <= #DLY 10'd0 ;
            in_dat_hld205[9:0] <= #DLY 10'd0 ;
            in_dat_hld206[9:0] <= #DLY 10'd0 ;
            in_dat_hld207[9:0] <= #DLY 10'd0 ;
            in_dat_hld208[9:0] <= #DLY 10'd0 ;
            in_dat_hld209[9:0] <= #DLY 10'd0 ;
            in_dat_hld210[9:0] <= #DLY 10'd0 ;
            in_dat_hld211[9:0] <= #DLY 10'd0 ;
            in_dat_hld212[9:0] <= #DLY 10'd0 ;
            in_dat_hld213[9:0] <= #DLY 10'd0 ;
            in_dat_hld214[9:0] <= #DLY 10'd0 ;
            in_dat_hld215[9:0] <= #DLY 10'd0 ;
            in_dat_hld216[9:0] <= #DLY 10'd0 ;
            in_dat_hld217[9:0] <= #DLY 10'd0 ;
            in_dat_hld218[9:0] <= #DLY 10'd0 ;
            in_dat_hld219[9:0] <= #DLY 10'd0 ;
            in_dat_hld220[9:0] <= #DLY 10'd0 ;
            in_dat_hld221[9:0] <= #DLY 10'd0 ;
            in_dat_hld222[9:0] <= #DLY 10'd0 ;
            in_dat_hld223[9:0] <= #DLY 10'd0 ;
            in_dat_hld224[9:0] <= #DLY 10'd0 ;
            in_dat_hld225[9:0] <= #DLY 10'd0 ;
            in_dat_hld226[9:0] <= #DLY 10'd0 ;
            in_dat_hld227[9:0] <= #DLY 10'd0 ;
            in_dat_hld228[9:0] <= #DLY 10'd0 ;
            in_dat_hld229[9:0] <= #DLY 10'd0 ;
            in_dat_hld230[9:0] <= #DLY 10'd0 ;
            in_dat_hld231[9:0] <= #DLY 10'd0 ;
            in_dat_hld232[9:0] <= #DLY 10'd0 ;
            in_dat_hld233[9:0] <= #DLY 10'd0 ;
            in_dat_hld234[9:0] <= #DLY 10'd0 ;
            in_dat_hld235[9:0] <= #DLY 10'd0 ;
            in_dat_hld236[9:0] <= #DLY 10'd0 ;
            in_dat_hld237[9:0] <= #DLY 10'd0 ;
            in_dat_hld238[9:0] <= #DLY 10'd0 ;
            in_dat_hld239[9:0] <= #DLY 10'd0 ;
            in_dat_hld240[9:0] <= #DLY 10'd0 ;
            in_dat_hld241[9:0] <= #DLY 10'd0 ;
            in_dat_hld242[9:0] <= #DLY 10'd0 ;
            in_dat_hld243[9:0] <= #DLY 10'd0 ;
            in_dat_hld244[9:0] <= #DLY 10'd0 ;
            in_dat_hld245[9:0] <= #DLY 10'd0 ;
            in_dat_hld246[9:0] <= #DLY 10'd0 ;
            in_dat_hld247[9:0] <= #DLY 10'd0 ;
            in_dat_hld248[9:0] <= #DLY 10'd0 ;
            in_dat_hld249[9:0] <= #DLY 10'd0 ;
            in_dat_hld250[9:0] <= #DLY 10'd0 ;
            in_dat_hld251[9:0] <= #DLY 10'd0 ;
            in_dat_hld252[9:0] <= #DLY 10'd0 ;
            in_dat_hld253[9:0] <= #DLY 10'd0 ;
            in_dat_hld254[9:0] <= #DLY 10'd0 ;
            in_dat_hld255[9:0] <= #DLY 10'd0 ;
            in_dat_hld256[9:0] <= #DLY 10'd0 ;
            in_dat_hld257[9:0] <= #DLY 10'd0 ;
            in_dat_hld258[9:0] <= #DLY 10'd0 ;
            in_dat_hld259[9:0] <= #DLY 10'd0 ;
            in_dat_hld260[9:0] <= #DLY 10'd0 ;
            in_dat_hld261[9:0] <= #DLY 10'd0 ;
            in_dat_hld262[9:0] <= #DLY 10'd0 ;
            in_dat_hld263[9:0] <= #DLY 10'd0 ;
            in_dat_hld264[9:0] <= #DLY 10'd0 ;
            in_dat_hld265[9:0] <= #DLY 10'd0 ;
            in_dat_hld266[9:0] <= #DLY 10'd0 ;
            in_dat_hld267[9:0] <= #DLY 10'd0 ;
            in_dat_hld268[9:0] <= #DLY 10'd0 ;
            in_dat_hld269[9:0] <= #DLY 10'd0 ;
            in_dat_hld270[9:0] <= #DLY 10'd0 ;
            in_dat_hld271[9:0] <= #DLY 10'd0 ;
            in_dat_hld272[9:0] <= #DLY 10'd0 ;
            in_dat_hld273[9:0] <= #DLY 10'd0 ;
            in_dat_hld274[9:0] <= #DLY 10'd0 ;
            in_dat_hld275[9:0] <= #DLY 10'd0 ;
            in_dat_hld276[9:0] <= #DLY 10'd0 ;
            in_dat_hld277[9:0] <= #DLY 10'd0 ;
            in_dat_hld278[9:0] <= #DLY 10'd0 ;
            in_dat_hld279[9:0] <= #DLY 10'd0 ;
            in_dat_hld280[9:0] <= #DLY 10'd0 ;
            in_dat_hld281[9:0] <= #DLY 10'd0 ;
            in_dat_hld282[9:0] <= #DLY 10'd0 ;
            in_dat_hld283[9:0] <= #DLY 10'd0 ;
            in_dat_hld284[9:0] <= #DLY 10'd0 ;
            in_dat_hld285[9:0] <= #DLY 10'd0 ;
            in_dat_hld286[9:0] <= #DLY 10'd0 ;
            in_dat_hld287[9:0] <= #DLY 10'd0 ;
            in_dat_hld288[9:0] <= #DLY 10'd0 ;
            in_dat_hld289[9:0] <= #DLY 10'd0 ;
            in_dat_hld290[9:0] <= #DLY 10'd0 ;
            in_dat_hld291[9:0] <= #DLY 10'd0 ;
            in_dat_hld292[9:0] <= #DLY 10'd0 ;
            in_dat_hld293[9:0] <= #DLY 10'd0 ;
            in_dat_hld294[9:0] <= #DLY 10'd0 ;
            in_dat_hld295[9:0] <= #DLY 10'd0 ;
            in_dat_hld296[9:0] <= #DLY 10'd0 ;
            in_dat_hld297[9:0] <= #DLY 10'd0 ;
            in_dat_hld298[9:0] <= #DLY 10'd0 ;
            in_dat_hld299[9:0] <= #DLY 10'd0 ;
            in_dat_hld300[9:0] <= #DLY 10'd0 ;
            in_dat_hld301[9:0] <= #DLY 10'd0 ;
            in_dat_hld302[9:0] <= #DLY 10'd0 ;
            in_dat_hld303[9:0] <= #DLY 10'd0 ;
            in_dat_hld304[9:0] <= #DLY 10'd0 ;
            in_dat_hld305[9:0] <= #DLY 10'd0 ;
            in_dat_hld306[9:0] <= #DLY 10'd0 ;
            in_dat_hld307[9:0] <= #DLY 10'd0 ;
            in_dat_hld308[9:0] <= #DLY 10'd0 ;
            in_dat_hld309[9:0] <= #DLY 10'd0 ;
            in_dat_hld310[9:0] <= #DLY 10'd0 ;
            in_dat_hld311[9:0] <= #DLY 10'd0 ;
            in_dat_hld312[9:0] <= #DLY 10'd0 ;
            in_dat_hld313[9:0] <= #DLY 10'd0 ;
            in_dat_hld314[9:0] <= #DLY 10'd0 ;
            in_dat_hld315[9:0] <= #DLY 10'd0 ;
            in_dat_hld316[9:0] <= #DLY 10'd0 ;
            in_dat_hld317[9:0] <= #DLY 10'd0 ;
            in_dat_hld318[9:0] <= #DLY 10'd0 ;
            in_dat_hld319[9:0] <= #DLY 10'd0 ;
            in_dat_hld320[9:0] <= #DLY 10'd0 ;
            in_dat_hld321[9:0] <= #DLY 10'd0 ;
            in_dat_hld322[9:0] <= #DLY 10'd0 ;
            in_dat_hld323[9:0] <= #DLY 10'd0 ;
            in_dat_hld324[9:0] <= #DLY 10'd0 ;
            in_dat_hld325[9:0] <= #DLY 10'd0 ;
            in_dat_hld326[9:0] <= #DLY 10'd0 ;
            in_dat_hld327[9:0] <= #DLY 10'd0 ;
            in_dat_hld328[9:0] <= #DLY 10'd0 ;
            in_dat_hld329[9:0] <= #DLY 10'd0 ;
            in_dat_hld330[9:0] <= #DLY 10'd0 ;
            in_dat_hld331[9:0] <= #DLY 10'd0 ;
            in_dat_hld332[9:0] <= #DLY 10'd0 ;
            in_dat_hld333[9:0] <= #DLY 10'd0 ;
            in_dat_hld334[9:0] <= #DLY 10'd0 ;
            in_dat_hld335[9:0] <= #DLY 10'd0 ;
            in_dat_hld336[9:0] <= #DLY 10'd0 ;
            in_dat_hld337[9:0] <= #DLY 10'd0 ;
            in_dat_hld338[9:0] <= #DLY 10'd0 ;
            in_dat_hld339[9:0] <= #DLY 10'd0 ;
            in_dat_hld340[9:0] <= #DLY 10'd0 ;
            in_dat_hld341[9:0] <= #DLY 10'd0 ;
            in_dat_hld342[9:0] <= #DLY 10'd0 ;
            in_dat_hld343[9:0] <= #DLY 10'd0 ;
            in_dat_hld344[9:0] <= #DLY 10'd0 ;
            in_dat_hld345[9:0] <= #DLY 10'd0 ;
            in_dat_hld346[9:0] <= #DLY 10'd0 ;
            in_dat_hld347[9:0] <= #DLY 10'd0 ;
            in_dat_hld348[9:0] <= #DLY 10'd0 ;
            in_dat_hld349[9:0] <= #DLY 10'd0 ;
            in_dat_hld350[9:0] <= #DLY 10'd0 ;
            in_dat_hld351[9:0] <= #DLY 10'd0 ;
            in_dat_hld352[9:0] <= #DLY 10'd0 ;
            in_dat_hld353[9:0] <= #DLY 10'd0 ;
            in_dat_hld354[9:0] <= #DLY 10'd0 ;
            in_dat_hld355[9:0] <= #DLY 10'd0 ;
            in_dat_hld356[9:0] <= #DLY 10'd0 ;
            in_dat_hld357[9:0] <= #DLY 10'd0 ;
            in_dat_hld358[9:0] <= #DLY 10'd0 ;
            in_dat_hld359[9:0] <= #DLY 10'd0 ;
            in_dat_hld360[9:0] <= #DLY 10'd0 ;
            in_dat_hld361[9:0] <= #DLY 10'd0 ;
            in_dat_hld362[9:0] <= #DLY 10'd0 ;
            in_dat_hld363[9:0] <= #DLY 10'd0 ;
            in_dat_hld364[9:0] <= #DLY 10'd0 ;
            in_dat_hld365[9:0] <= #DLY 10'd0 ;
            in_dat_hld366[9:0] <= #DLY 10'd0 ;
            in_dat_hld367[9:0] <= #DLY 10'd0 ;
            in_dat_hld368[9:0] <= #DLY 10'd0 ;
            in_dat_hld369[9:0] <= #DLY 10'd0 ;
            in_dat_hld370[9:0] <= #DLY 10'd0 ;
            in_dat_hld371[9:0] <= #DLY 10'd0 ;
            in_dat_hld372[9:0] <= #DLY 10'd0 ;
            in_dat_hld373[9:0] <= #DLY 10'd0 ;
            in_dat_hld374[9:0] <= #DLY 10'd0 ;
            in_dat_hld375[9:0] <= #DLY 10'd0 ;
            in_dat_hld376[9:0] <= #DLY 10'd0 ;
            in_dat_hld377[9:0] <= #DLY 10'd0 ;
            in_dat_hld378[9:0] <= #DLY 10'd0 ;
            in_dat_hld379[9:0] <= #DLY 10'd0 ;
            in_dat_hld380[9:0] <= #DLY 10'd0 ;
            in_dat_hld381[9:0] <= #DLY 10'd0 ;
            in_dat_hld382[9:0] <= #DLY 10'd0 ;
            in_dat_hld383[9:0] <= #DLY 10'd0 ;
            in_dat_hld384[9:0] <= #DLY 10'd0 ;
            in_dat_hld385[9:0] <= #DLY 10'd0 ;
            in_dat_hld386[9:0] <= #DLY 10'd0 ;
            in_dat_hld387[9:0] <= #DLY 10'd0 ;
            in_dat_hld388[9:0] <= #DLY 10'd0 ;
            in_dat_hld389[9:0] <= #DLY 10'd0 ;
            in_dat_hld390[9:0] <= #DLY 10'd0 ;
            in_dat_hld391[9:0] <= #DLY 10'd0 ;
            in_dat_hld392[9:0] <= #DLY 10'd0 ;
            in_dat_hld393[9:0] <= #DLY 10'd0 ;
            in_dat_hld394[9:0] <= #DLY 10'd0 ;
            in_dat_hld395[9:0] <= #DLY 10'd0 ;
            in_dat_hld396[9:0] <= #DLY 10'd0 ;
            in_dat_hld397[9:0] <= #DLY 10'd0 ;
            in_dat_hld398[9:0] <= #DLY 10'd0 ;
            in_dat_hld399[9:0] <= #DLY 10'd0 ;
            in_dat_hld400[9:0] <= #DLY 10'd0 ;
            in_dat_hld401[9:0] <= #DLY 10'd0 ;
            in_dat_hld402[9:0] <= #DLY 10'd0 ;
            in_dat_hld403[9:0] <= #DLY 10'd0 ;
            in_dat_hld404[9:0] <= #DLY 10'd0 ;
            in_dat_hld405[9:0] <= #DLY 10'd0 ;
            in_dat_hld406[9:0] <= #DLY 10'd0 ;
            in_dat_hld407[9:0] <= #DLY 10'd0 ;
            in_dat_hld408[9:0] <= #DLY 10'd0 ;
            in_dat_hld409[9:0] <= #DLY 10'd0 ;
            in_dat_hld410[9:0] <= #DLY 10'd0 ;
            in_dat_hld411[9:0] <= #DLY 10'd0 ;
            in_dat_hld412[9:0] <= #DLY 10'd0 ;
            in_dat_hld413[9:0] <= #DLY 10'd0 ;
            in_dat_hld414[9:0] <= #DLY 10'd0 ;
            in_dat_hld415[9:0] <= #DLY 10'd0 ;
            in_dat_hld416[9:0] <= #DLY 10'd0 ;
            in_dat_hld417[9:0] <= #DLY 10'd0 ;
            in_dat_hld418[9:0] <= #DLY 10'd0 ;
            in_dat_hld419[9:0] <= #DLY 10'd0 ;
            in_dat_hld420[9:0] <= #DLY 10'd0 ;
            in_dat_hld421[9:0] <= #DLY 10'd0 ;
            in_dat_hld422[9:0] <= #DLY 10'd0 ;
            in_dat_hld423[9:0] <= #DLY 10'd0 ;
            in_dat_hld424[9:0] <= #DLY 10'd0 ;
            in_dat_hld425[9:0] <= #DLY 10'd0 ;
            in_dat_hld426[9:0] <= #DLY 10'd0 ;
            in_dat_hld427[9:0] <= #DLY 10'd0 ;
            in_dat_hld428[9:0] <= #DLY 10'd0 ;
            in_dat_hld429[9:0] <= #DLY 10'd0 ;
            in_dat_hld430[9:0] <= #DLY 10'd0 ;
            in_dat_hld431[9:0] <= #DLY 10'd0 ;
            in_dat_hld432[9:0] <= #DLY 10'd0 ;
            in_dat_hld433[9:0] <= #DLY 10'd0 ;
            in_dat_hld434[9:0] <= #DLY 10'd0 ;
            in_dat_hld435[9:0] <= #DLY 10'd0 ;
            in_dat_hld436[9:0] <= #DLY 10'd0 ;
            in_dat_hld437[9:0] <= #DLY 10'd0 ;
            in_dat_hld438[9:0] <= #DLY 10'd0 ;
            in_dat_hld439[9:0] <= #DLY 10'd0 ;
            in_dat_hld440[9:0] <= #DLY 10'd0 ;
            in_dat_hld441[9:0] <= #DLY 10'd0 ;
            in_dat_hld442[9:0] <= #DLY 10'd0 ;
            in_dat_hld443[9:0] <= #DLY 10'd0 ;
            in_dat_hld444[9:0] <= #DLY 10'd0 ;
            in_dat_hld445[9:0] <= #DLY 10'd0 ;
            in_dat_hld446[9:0] <= #DLY 10'd0 ;
            in_dat_hld447[9:0] <= #DLY 10'd0 ;
            in_dat_hld448[9:0] <= #DLY 10'd0 ;
            in_dat_hld449[9:0] <= #DLY 10'd0 ;
            in_dat_hld450[9:0] <= #DLY 10'd0 ;
            in_dat_hld451[9:0] <= #DLY 10'd0 ;
            in_dat_hld452[9:0] <= #DLY 10'd0 ;
            in_dat_hld453[9:0] <= #DLY 10'd0 ;
            in_dat_hld454[9:0] <= #DLY 10'd0 ;
            in_dat_hld455[9:0] <= #DLY 10'd0 ;
            in_dat_hld456[9:0] <= #DLY 10'd0 ;
            in_dat_hld457[9:0] <= #DLY 10'd0 ;
            in_dat_hld458[9:0] <= #DLY 10'd0 ;
            in_dat_hld459[9:0] <= #DLY 10'd0 ;
            in_dat_hld460[9:0] <= #DLY 10'd0 ;
            in_dat_hld461[9:0] <= #DLY 10'd0 ;
            in_dat_hld462[9:0] <= #DLY 10'd0 ;
            in_dat_hld463[9:0] <= #DLY 10'd0 ;
            in_dat_hld464[9:0] <= #DLY 10'd0 ;
            in_dat_hld465[9:0] <= #DLY 10'd0 ;
            in_dat_hld466[9:0] <= #DLY 10'd0 ;
            in_dat_hld467[9:0] <= #DLY 10'd0 ;
            in_dat_hld468[9:0] <= #DLY 10'd0 ;
            in_dat_hld469[9:0] <= #DLY 10'd0 ;
            in_dat_hld470[9:0] <= #DLY 10'd0 ;
            in_dat_hld471[9:0] <= #DLY 10'd0 ;
            in_dat_hld472[9:0] <= #DLY 10'd0 ;
            in_dat_hld473[9:0] <= #DLY 10'd0 ;
            in_dat_hld474[9:0] <= #DLY 10'd0 ;
            in_dat_hld475[9:0] <= #DLY 10'd0 ;
            in_dat_hld476[9:0] <= #DLY 10'd0 ;
            in_dat_hld477[9:0] <= #DLY 10'd0 ;
            in_dat_hld478[9:0] <= #DLY 10'd0 ;
            in_dat_hld479[9:0] <= #DLY 10'd0 ;
            in_dat_hld480[9:0] <= #DLY 10'd0 ;
            in_dat_hld481[9:0] <= #DLY 10'd0 ;
            in_dat_hld482[9:0] <= #DLY 10'd0 ;
            in_dat_hld483[9:0] <= #DLY 10'd0 ;
            in_dat_hld484[9:0] <= #DLY 10'd0 ;
            in_dat_hld485[9:0] <= #DLY 10'd0 ;
            in_dat_hld486[9:0] <= #DLY 10'd0 ;
            in_dat_hld487[9:0] <= #DLY 10'd0 ;
            in_dat_hld488[9:0] <= #DLY 10'd0 ;
            in_dat_hld489[9:0] <= #DLY 10'd0 ;
            in_dat_hld490[9:0] <= #DLY 10'd0 ;
            in_dat_hld491[9:0] <= #DLY 10'd0 ;
            in_dat_hld492[9:0] <= #DLY 10'd0 ;
            in_dat_hld493[9:0] <= #DLY 10'd0 ;
            in_dat_hld494[9:0] <= #DLY 10'd0 ;
            in_dat_hld495[9:0] <= #DLY 10'd0 ;
            in_dat_hld496[9:0] <= #DLY 10'd0 ;
            in_dat_hld497[9:0] <= #DLY 10'd0 ;
            in_dat_hld498[9:0] <= #DLY 10'd0 ;
            in_dat_hld499[9:0] <= #DLY 10'd0 ;
            in_dat_hld500[9:0] <= #DLY 10'd0 ;
            in_dat_hld501[9:0] <= #DLY 10'd0 ;
            in_dat_hld502[9:0] <= #DLY 10'd0 ;
            in_dat_hld503[9:0] <= #DLY 10'd0 ;
            in_dat_hld504[9:0] <= #DLY 10'd0 ;
            in_dat_hld505[9:0] <= #DLY 10'd0 ;
            in_dat_hld506[9:0] <= #DLY 10'd0 ;
            in_dat_hld507[9:0] <= #DLY 10'd0 ;
            in_dat_hld508[9:0] <= #DLY 10'd0 ;
            in_dat_hld509[9:0] <= #DLY 10'd0 ;
            in_dat_hld510[9:0] <= #DLY 10'd0 ;
            in_dat_hld511[9:0] <= #DLY 10'd0 ;
            in_dat_hld512[9:0] <= #DLY 10'd0 ;
		end else begin
		    if(pipeline_cnt[32] & (cyc32_cnt_dd1[5:0]==6'd31)) begin
                in_dat_hld01[9:0]  <= #DLY in_dat_wire01[9:0]  ;
                in_dat_hld02[9:0]  <= #DLY in_dat_wire02[9:0]  ;
                in_dat_hld03[9:0]  <= #DLY in_dat_wire03[9:0]  ;
                in_dat_hld04[9:0]  <= #DLY in_dat_wire04[9:0]  ;
                in_dat_hld05[9:0]  <= #DLY in_dat_wire05[9:0]  ;
                in_dat_hld06[9:0]  <= #DLY in_dat_wire06[9:0]  ;
                in_dat_hld07[9:0]  <= #DLY in_dat_wire07[9:0]  ;
                in_dat_hld08[9:0]  <= #DLY in_dat_wire08[9:0]  ;
                in_dat_hld09[9:0]  <= #DLY in_dat_wire09[9:0]  ;
                in_dat_hld10[9:0]  <= #DLY in_dat_wire10[9:0]  ;
                in_dat_hld11[9:0]  <= #DLY in_dat_wire11[9:0]  ;
                in_dat_hld12[9:0]  <= #DLY in_dat_wire12[9:0]  ;
                in_dat_hld13[9:0]  <= #DLY in_dat_wire13[9:0]  ;
                in_dat_hld14[9:0]  <= #DLY in_dat_wire14[9:0]  ;
                in_dat_hld15[9:0]  <= #DLY in_dat_wire15[9:0]  ;
                in_dat_hld16[9:0]  <= #DLY in_dat_wire16[9:0]  ;
                in_dat_hld17[9:0]  <= #DLY in_dat_wire17[9:0]  ;
                in_dat_hld18[9:0]  <= #DLY in_dat_wire18[9:0]  ;
                in_dat_hld19[9:0]  <= #DLY in_dat_wire19[9:0]  ;
                in_dat_hld20[9:0]  <= #DLY in_dat_wire20[9:0]  ;
                in_dat_hld21[9:0]  <= #DLY in_dat_wire21[9:0]  ;
                in_dat_hld22[9:0]  <= #DLY in_dat_wire22[9:0]  ;
                in_dat_hld23[9:0]  <= #DLY in_dat_wire23[9:0]  ;
                in_dat_hld24[9:0]  <= #DLY in_dat_wire24[9:0]  ;
                in_dat_hld25[9:0]  <= #DLY in_dat_wire25[9:0]  ;
                in_dat_hld26[9:0]  <= #DLY in_dat_wire26[9:0]  ;
                in_dat_hld27[9:0]  <= #DLY in_dat_wire27[9:0]  ;
                in_dat_hld28[9:0]  <= #DLY in_dat_wire28[9:0]  ;
                in_dat_hld29[9:0]  <= #DLY in_dat_wire29[9:0]  ;
                in_dat_hld30[9:0]  <= #DLY in_dat_wire30[9:0]  ;
                in_dat_hld31[9:0]  <= #DLY in_dat_wire31[9:0]  ;
                in_dat_hld32[9:0]  <= #DLY in_dat_wire32[9:0]  ;
                in_dat_hld33[9:0]  <= #DLY in_dat_wire33[9:0]  ;
                in_dat_hld34[9:0]  <= #DLY in_dat_wire34[9:0]  ;
                in_dat_hld35[9:0]  <= #DLY in_dat_wire35[9:0]  ;
                in_dat_hld36[9:0]  <= #DLY in_dat_wire36[9:0]  ;
                in_dat_hld37[9:0]  <= #DLY in_dat_wire37[9:0]  ;
                in_dat_hld38[9:0]  <= #DLY in_dat_wire38[9:0]  ;
                in_dat_hld39[9:0]  <= #DLY in_dat_wire39[9:0]  ;
                in_dat_hld40[9:0]  <= #DLY in_dat_wire40[9:0]  ;
                in_dat_hld41[9:0]  <= #DLY in_dat_wire41[9:0]  ;
                in_dat_hld42[9:0]  <= #DLY in_dat_wire42[9:0]  ;
                in_dat_hld43[9:0]  <= #DLY in_dat_wire43[9:0]  ;
                in_dat_hld44[9:0]  <= #DLY in_dat_wire44[9:0]  ;
                in_dat_hld45[9:0]  <= #DLY in_dat_wire45[9:0]  ;
                in_dat_hld46[9:0]  <= #DLY in_dat_wire46[9:0]  ;
                in_dat_hld47[9:0]  <= #DLY in_dat_wire47[9:0]  ;
                in_dat_hld48[9:0]  <= #DLY in_dat_wire48[9:0]  ;
                in_dat_hld49[9:0]  <= #DLY in_dat_wire49[9:0]  ;
                in_dat_hld50[9:0]  <= #DLY in_dat_wire50[9:0]  ;
                in_dat_hld51[9:0]  <= #DLY in_dat_wire51[9:0]  ;
                in_dat_hld52[9:0]  <= #DLY in_dat_wire52[9:0]  ;
                in_dat_hld53[9:0]  <= #DLY in_dat_wire53[9:0]  ;
                in_dat_hld54[9:0]  <= #DLY in_dat_wire54[9:0]  ;
                in_dat_hld55[9:0]  <= #DLY in_dat_wire55[9:0]  ;
                in_dat_hld56[9:0]  <= #DLY in_dat_wire56[9:0]  ;
                in_dat_hld57[9:0]  <= #DLY in_dat_wire57[9:0]  ;
                in_dat_hld58[9:0]  <= #DLY in_dat_wire58[9:0]  ;
                in_dat_hld59[9:0]  <= #DLY in_dat_wire59[9:0]  ;
                in_dat_hld60[9:0]  <= #DLY in_dat_wire60[9:0]  ;
                in_dat_hld61[9:0]  <= #DLY in_dat_wire61[9:0]  ;
                in_dat_hld62[9:0]  <= #DLY in_dat_wire62[9:0]  ;
                in_dat_hld63[9:0]  <= #DLY in_dat_wire63[9:0]  ;
                in_dat_hld64[9:0]  <= #DLY in_dat_wire64[9:0]  ;
                in_dat_hld65[9:0]  <= #DLY in_dat_wire65[9:0]  ;
                in_dat_hld66[9:0]  <= #DLY in_dat_wire66[9:0]  ;
                in_dat_hld67[9:0]  <= #DLY in_dat_wire67[9:0]  ;
                in_dat_hld68[9:0]  <= #DLY in_dat_wire68[9:0]  ;
                in_dat_hld69[9:0]  <= #DLY in_dat_wire69[9:0]  ;
                in_dat_hld70[9:0]  <= #DLY in_dat_wire70[9:0]  ;
                in_dat_hld71[9:0]  <= #DLY in_dat_wire71[9:0]  ;
                in_dat_hld72[9:0]  <= #DLY in_dat_wire72[9:0]  ;
                in_dat_hld73[9:0]  <= #DLY in_dat_wire73[9:0]  ;
                in_dat_hld74[9:0]  <= #DLY in_dat_wire74[9:0]  ;
                in_dat_hld75[9:0]  <= #DLY in_dat_wire75[9:0]  ;
                in_dat_hld76[9:0]  <= #DLY in_dat_wire76[9:0]  ;
                in_dat_hld77[9:0]  <= #DLY in_dat_wire77[9:0]  ;
                in_dat_hld78[9:0]  <= #DLY in_dat_wire78[9:0]  ;
                in_dat_hld79[9:0]  <= #DLY in_dat_wire79[9:0]  ;
                in_dat_hld80[9:0]  <= #DLY in_dat_wire80[9:0]  ;
                in_dat_hld81[9:0]  <= #DLY in_dat_wire81[9:0]  ;
                in_dat_hld82[9:0]  <= #DLY in_dat_wire82[9:0]  ;
                in_dat_hld83[9:0]  <= #DLY in_dat_wire83[9:0]  ;
                in_dat_hld84[9:0]  <= #DLY in_dat_wire84[9:0]  ;
                in_dat_hld85[9:0]  <= #DLY in_dat_wire85[9:0]  ;
                in_dat_hld86[9:0]  <= #DLY in_dat_wire86[9:0]  ;
                in_dat_hld87[9:0]  <= #DLY in_dat_wire87[9:0]  ;
                in_dat_hld88[9:0]  <= #DLY in_dat_wire88[9:0]  ;
                in_dat_hld89[9:0]  <= #DLY in_dat_wire89[9:0]  ;
                in_dat_hld90[9:0]  <= #DLY in_dat_wire90[9:0]  ;
                in_dat_hld91[9:0]  <= #DLY in_dat_wire91[9:0]  ;
                in_dat_hld92[9:0]  <= #DLY in_dat_wire92[9:0]  ;
                in_dat_hld93[9:0]  <= #DLY in_dat_wire93[9:0]  ;
                in_dat_hld94[9:0]  <= #DLY in_dat_wire94[9:0]  ;
                in_dat_hld95[9:0]  <= #DLY in_dat_wire95[9:0]  ;
                in_dat_hld96[9:0]  <= #DLY in_dat_wire96[9:0]  ;
                in_dat_hld97[9:0]  <= #DLY in_dat_wire97[9:0]  ;
                in_dat_hld98[9:0]  <= #DLY in_dat_wire98[9:0]  ;
                in_dat_hld99[9:0]  <= #DLY in_dat_wire99[9:0]  ;
                in_dat_hld100[9:0] <= #DLY in_dat_wire100[9:0] ;
                in_dat_hld101[9:0] <= #DLY in_dat_wire101[9:0] ;
                in_dat_hld102[9:0] <= #DLY in_dat_wire102[9:0] ;
                in_dat_hld103[9:0] <= #DLY in_dat_wire103[9:0] ;
                in_dat_hld104[9:0] <= #DLY in_dat_wire104[9:0] ;
                in_dat_hld105[9:0] <= #DLY in_dat_wire105[9:0] ;
                in_dat_hld106[9:0] <= #DLY in_dat_wire106[9:0] ;
                in_dat_hld107[9:0] <= #DLY in_dat_wire107[9:0] ;
                in_dat_hld108[9:0] <= #DLY in_dat_wire108[9:0] ;
                in_dat_hld109[9:0] <= #DLY in_dat_wire109[9:0] ;
                in_dat_hld110[9:0] <= #DLY in_dat_wire110[9:0] ;
                in_dat_hld111[9:0] <= #DLY in_dat_wire111[9:0] ;
                in_dat_hld112[9:0] <= #DLY in_dat_wire112[9:0] ;
                in_dat_hld113[9:0] <= #DLY in_dat_wire113[9:0] ;
                in_dat_hld114[9:0] <= #DLY in_dat_wire114[9:0] ;
                in_dat_hld115[9:0] <= #DLY in_dat_wire115[9:0] ;
                in_dat_hld116[9:0] <= #DLY in_dat_wire116[9:0] ;
                in_dat_hld117[9:0] <= #DLY in_dat_wire117[9:0] ;
                in_dat_hld118[9:0] <= #DLY in_dat_wire118[9:0] ;
                in_dat_hld119[9:0] <= #DLY in_dat_wire119[9:0] ;
                in_dat_hld120[9:0] <= #DLY in_dat_wire120[9:0] ;
                in_dat_hld121[9:0] <= #DLY in_dat_wire121[9:0] ;
                in_dat_hld122[9:0] <= #DLY in_dat_wire122[9:0] ;
                in_dat_hld123[9:0] <= #DLY in_dat_wire123[9:0] ;
                in_dat_hld124[9:0] <= #DLY in_dat_wire124[9:0] ;
                in_dat_hld125[9:0] <= #DLY in_dat_wire125[9:0] ;
                in_dat_hld126[9:0] <= #DLY in_dat_wire126[9:0] ;
                in_dat_hld127[9:0] <= #DLY in_dat_wire127[9:0] ;
                in_dat_hld128[9:0] <= #DLY in_dat_wire128[9:0] ;
                in_dat_hld129[9:0] <= #DLY in_dat_wire129[9:0] ;
                in_dat_hld130[9:0] <= #DLY in_dat_wire130[9:0] ;
                in_dat_hld131[9:0] <= #DLY in_dat_wire131[9:0] ;
                in_dat_hld132[9:0] <= #DLY in_dat_wire132[9:0] ;
                in_dat_hld133[9:0] <= #DLY in_dat_wire133[9:0] ;
                in_dat_hld134[9:0] <= #DLY in_dat_wire134[9:0] ;
                in_dat_hld135[9:0] <= #DLY in_dat_wire135[9:0] ;
                in_dat_hld136[9:0] <= #DLY in_dat_wire136[9:0] ;
                in_dat_hld137[9:0] <= #DLY in_dat_wire137[9:0] ;
                in_dat_hld138[9:0] <= #DLY in_dat_wire138[9:0] ;
                in_dat_hld139[9:0] <= #DLY in_dat_wire139[9:0] ;
                in_dat_hld140[9:0] <= #DLY in_dat_wire140[9:0] ;
                in_dat_hld141[9:0] <= #DLY in_dat_wire141[9:0] ;
                in_dat_hld142[9:0] <= #DLY in_dat_wire142[9:0] ;
                in_dat_hld143[9:0] <= #DLY in_dat_wire143[9:0] ;
                in_dat_hld144[9:0] <= #DLY in_dat_wire144[9:0] ;
                in_dat_hld145[9:0] <= #DLY in_dat_wire145[9:0] ;
                in_dat_hld146[9:0] <= #DLY in_dat_wire146[9:0] ;
                in_dat_hld147[9:0] <= #DLY in_dat_wire147[9:0] ;
                in_dat_hld148[9:0] <= #DLY in_dat_wire148[9:0] ;
                in_dat_hld149[9:0] <= #DLY in_dat_wire149[9:0] ;
                in_dat_hld150[9:0] <= #DLY in_dat_wire150[9:0] ;
                in_dat_hld151[9:0] <= #DLY in_dat_wire151[9:0] ;
                in_dat_hld152[9:0] <= #DLY in_dat_wire152[9:0] ;
                in_dat_hld153[9:0] <= #DLY in_dat_wire153[9:0] ;
                in_dat_hld154[9:0] <= #DLY in_dat_wire154[9:0] ;
                in_dat_hld155[9:0] <= #DLY in_dat_wire155[9:0] ;
                in_dat_hld156[9:0] <= #DLY in_dat_wire156[9:0] ;
                in_dat_hld157[9:0] <= #DLY in_dat_wire157[9:0] ;
                in_dat_hld158[9:0] <= #DLY in_dat_wire158[9:0] ;
                in_dat_hld159[9:0] <= #DLY in_dat_wire159[9:0] ;
                in_dat_hld160[9:0] <= #DLY in_dat_wire160[9:0] ;
                in_dat_hld161[9:0] <= #DLY in_dat_wire161[9:0] ;
                in_dat_hld162[9:0] <= #DLY in_dat_wire162[9:0] ;
                in_dat_hld163[9:0] <= #DLY in_dat_wire163[9:0] ;
                in_dat_hld164[9:0] <= #DLY in_dat_wire164[9:0] ;
                in_dat_hld165[9:0] <= #DLY in_dat_wire165[9:0] ;
                in_dat_hld166[9:0] <= #DLY in_dat_wire166[9:0] ;
                in_dat_hld167[9:0] <= #DLY in_dat_wire167[9:0] ;
                in_dat_hld168[9:0] <= #DLY in_dat_wire168[9:0] ;
                in_dat_hld169[9:0] <= #DLY in_dat_wire169[9:0] ;
                in_dat_hld170[9:0] <= #DLY in_dat_wire170[9:0] ;
                in_dat_hld171[9:0] <= #DLY in_dat_wire171[9:0] ;
                in_dat_hld172[9:0] <= #DLY in_dat_wire172[9:0] ;
                in_dat_hld173[9:0] <= #DLY in_dat_wire173[9:0] ;
                in_dat_hld174[9:0] <= #DLY in_dat_wire174[9:0] ;
                in_dat_hld175[9:0] <= #DLY in_dat_wire175[9:0] ;
                in_dat_hld176[9:0] <= #DLY in_dat_wire176[9:0] ;
                in_dat_hld177[9:0] <= #DLY in_dat_wire177[9:0] ;
                in_dat_hld178[9:0] <= #DLY in_dat_wire178[9:0] ;
                in_dat_hld179[9:0] <= #DLY in_dat_wire179[9:0] ;
                in_dat_hld180[9:0] <= #DLY in_dat_wire180[9:0] ;
                in_dat_hld181[9:0] <= #DLY in_dat_wire181[9:0] ;
                in_dat_hld182[9:0] <= #DLY in_dat_wire182[9:0] ;
                in_dat_hld183[9:0] <= #DLY in_dat_wire183[9:0] ;
                in_dat_hld184[9:0] <= #DLY in_dat_wire184[9:0] ;
                in_dat_hld185[9:0] <= #DLY in_dat_wire185[9:0] ;
                in_dat_hld186[9:0] <= #DLY in_dat_wire186[9:0] ;
                in_dat_hld187[9:0] <= #DLY in_dat_wire187[9:0] ;
                in_dat_hld188[9:0] <= #DLY in_dat_wire188[9:0] ;
                in_dat_hld189[9:0] <= #DLY in_dat_wire189[9:0] ;
                in_dat_hld190[9:0] <= #DLY in_dat_wire190[9:0] ;
                in_dat_hld191[9:0] <= #DLY in_dat_wire191[9:0] ;
                in_dat_hld192[9:0] <= #DLY in_dat_wire192[9:0] ;
                in_dat_hld193[9:0] <= #DLY in_dat_wire193[9:0] ;
                in_dat_hld194[9:0] <= #DLY in_dat_wire194[9:0] ;
                in_dat_hld195[9:0] <= #DLY in_dat_wire195[9:0] ;
                in_dat_hld196[9:0] <= #DLY in_dat_wire196[9:0] ;
                in_dat_hld197[9:0] <= #DLY in_dat_wire197[9:0] ;
                in_dat_hld198[9:0] <= #DLY in_dat_wire198[9:0] ;
                in_dat_hld199[9:0] <= #DLY in_dat_wire199[9:0] ;
                in_dat_hld200[9:0] <= #DLY in_dat_wire200[9:0] ;
                in_dat_hld201[9:0] <= #DLY in_dat_wire201[9:0] ;
                in_dat_hld202[9:0] <= #DLY in_dat_wire202[9:0] ;
                in_dat_hld203[9:0] <= #DLY in_dat_wire203[9:0] ;
                in_dat_hld204[9:0] <= #DLY in_dat_wire204[9:0] ;
                in_dat_hld205[9:0] <= #DLY in_dat_wire205[9:0] ;
                in_dat_hld206[9:0] <= #DLY in_dat_wire206[9:0] ;
                in_dat_hld207[9:0] <= #DLY in_dat_wire207[9:0] ;
                in_dat_hld208[9:0] <= #DLY in_dat_wire208[9:0] ;
                in_dat_hld209[9:0] <= #DLY in_dat_wire209[9:0] ;
                in_dat_hld210[9:0] <= #DLY in_dat_wire210[9:0] ;
                in_dat_hld211[9:0] <= #DLY in_dat_wire211[9:0] ;
                in_dat_hld212[9:0] <= #DLY in_dat_wire212[9:0] ;
                in_dat_hld213[9:0] <= #DLY in_dat_wire213[9:0] ;
                in_dat_hld214[9:0] <= #DLY in_dat_wire214[9:0] ;
                in_dat_hld215[9:0] <= #DLY in_dat_wire215[9:0] ;
                in_dat_hld216[9:0] <= #DLY in_dat_wire216[9:0] ;
                in_dat_hld217[9:0] <= #DLY in_dat_wire217[9:0] ;
                in_dat_hld218[9:0] <= #DLY in_dat_wire218[9:0] ;
                in_dat_hld219[9:0] <= #DLY in_dat_wire219[9:0] ;
                in_dat_hld220[9:0] <= #DLY in_dat_wire220[9:0] ;
                in_dat_hld221[9:0] <= #DLY in_dat_wire221[9:0] ;
                in_dat_hld222[9:0] <= #DLY in_dat_wire222[9:0] ;
                in_dat_hld223[9:0] <= #DLY in_dat_wire223[9:0] ;
                in_dat_hld224[9:0] <= #DLY in_dat_wire224[9:0] ;
                in_dat_hld225[9:0] <= #DLY in_dat_wire225[9:0] ;
                in_dat_hld226[9:0] <= #DLY in_dat_wire226[9:0] ;
                in_dat_hld227[9:0] <= #DLY in_dat_wire227[9:0] ;
                in_dat_hld228[9:0] <= #DLY in_dat_wire228[9:0] ;
                in_dat_hld229[9:0] <= #DLY in_dat_wire229[9:0] ;
                in_dat_hld230[9:0] <= #DLY in_dat_wire230[9:0] ;
                in_dat_hld231[9:0] <= #DLY in_dat_wire231[9:0] ;
                in_dat_hld232[9:0] <= #DLY in_dat_wire232[9:0] ;
                in_dat_hld233[9:0] <= #DLY in_dat_wire233[9:0] ;
                in_dat_hld234[9:0] <= #DLY in_dat_wire234[9:0] ;
                in_dat_hld235[9:0] <= #DLY in_dat_wire235[9:0] ;
                in_dat_hld236[9:0] <= #DLY in_dat_wire236[9:0] ;
                in_dat_hld237[9:0] <= #DLY in_dat_wire237[9:0] ;
                in_dat_hld238[9:0] <= #DLY in_dat_wire238[9:0] ;
                in_dat_hld239[9:0] <= #DLY in_dat_wire239[9:0] ;
                in_dat_hld240[9:0] <= #DLY in_dat_wire240[9:0] ;
                in_dat_hld241[9:0] <= #DLY in_dat_wire241[9:0] ;
                in_dat_hld242[9:0] <= #DLY in_dat_wire242[9:0] ;
                in_dat_hld243[9:0] <= #DLY in_dat_wire243[9:0] ;
                in_dat_hld244[9:0] <= #DLY in_dat_wire244[9:0] ;
                in_dat_hld245[9:0] <= #DLY in_dat_wire245[9:0] ;
                in_dat_hld246[9:0] <= #DLY in_dat_wire246[9:0] ;
                in_dat_hld247[9:0] <= #DLY in_dat_wire247[9:0] ;
                in_dat_hld248[9:0] <= #DLY in_dat_wire248[9:0] ;
                in_dat_hld249[9:0] <= #DLY in_dat_wire249[9:0] ;
                in_dat_hld250[9:0] <= #DLY in_dat_wire250[9:0] ;
                in_dat_hld251[9:0] <= #DLY in_dat_wire251[9:0] ;
                in_dat_hld252[9:0] <= #DLY in_dat_wire252[9:0] ;
                in_dat_hld253[9:0] <= #DLY in_dat_wire253[9:0] ;
                in_dat_hld254[9:0] <= #DLY in_dat_wire254[9:0] ;
                in_dat_hld255[9:0] <= #DLY in_dat_wire255[9:0] ;
                in_dat_hld256[9:0] <= #DLY in_dat_wire256[9:0] ;
                in_dat_hld257[9:0] <= #DLY in_dat_wire257[9:0] ;
                in_dat_hld258[9:0] <= #DLY in_dat_wire258[9:0] ;
                in_dat_hld259[9:0] <= #DLY in_dat_wire259[9:0] ;
                in_dat_hld260[9:0] <= #DLY in_dat_wire260[9:0] ;
                in_dat_hld261[9:0] <= #DLY in_dat_wire261[9:0] ;
                in_dat_hld262[9:0] <= #DLY in_dat_wire262[9:0] ;
                in_dat_hld263[9:0] <= #DLY in_dat_wire263[9:0] ;
                in_dat_hld264[9:0] <= #DLY in_dat_wire264[9:0] ;
                in_dat_hld265[9:0] <= #DLY in_dat_wire265[9:0] ;
                in_dat_hld266[9:0] <= #DLY in_dat_wire266[9:0] ;
                in_dat_hld267[9:0] <= #DLY in_dat_wire267[9:0] ;
                in_dat_hld268[9:0] <= #DLY in_dat_wire268[9:0] ;
                in_dat_hld269[9:0] <= #DLY in_dat_wire269[9:0] ;
                in_dat_hld270[9:0] <= #DLY in_dat_wire270[9:0] ;
                in_dat_hld271[9:0] <= #DLY in_dat_wire271[9:0] ;
                in_dat_hld272[9:0] <= #DLY in_dat_wire272[9:0] ;
                in_dat_hld273[9:0] <= #DLY in_dat_wire273[9:0] ;
                in_dat_hld274[9:0] <= #DLY in_dat_wire274[9:0] ;
                in_dat_hld275[9:0] <= #DLY in_dat_wire275[9:0] ;
                in_dat_hld276[9:0] <= #DLY in_dat_wire276[9:0] ;
                in_dat_hld277[9:0] <= #DLY in_dat_wire277[9:0] ;
                in_dat_hld278[9:0] <= #DLY in_dat_wire278[9:0] ;
                in_dat_hld279[9:0] <= #DLY in_dat_wire279[9:0] ;
                in_dat_hld280[9:0] <= #DLY in_dat_wire280[9:0] ;
                in_dat_hld281[9:0] <= #DLY in_dat_wire281[9:0] ;
                in_dat_hld282[9:0] <= #DLY in_dat_wire282[9:0] ;
                in_dat_hld283[9:0] <= #DLY in_dat_wire283[9:0] ;
                in_dat_hld284[9:0] <= #DLY in_dat_wire284[9:0] ;
                in_dat_hld285[9:0] <= #DLY in_dat_wire285[9:0] ;
                in_dat_hld286[9:0] <= #DLY in_dat_wire286[9:0] ;
                in_dat_hld287[9:0] <= #DLY in_dat_wire287[9:0] ;
                in_dat_hld288[9:0] <= #DLY in_dat_wire288[9:0] ;
                in_dat_hld289[9:0] <= #DLY in_dat_wire289[9:0] ;
                in_dat_hld290[9:0] <= #DLY in_dat_wire290[9:0] ;
                in_dat_hld291[9:0] <= #DLY in_dat_wire291[9:0] ;
                in_dat_hld292[9:0] <= #DLY in_dat_wire292[9:0] ;
                in_dat_hld293[9:0] <= #DLY in_dat_wire293[9:0] ;
                in_dat_hld294[9:0] <= #DLY in_dat_wire294[9:0] ;
                in_dat_hld295[9:0] <= #DLY in_dat_wire295[9:0] ;
                in_dat_hld296[9:0] <= #DLY in_dat_wire296[9:0] ;
                in_dat_hld297[9:0] <= #DLY in_dat_wire297[9:0] ;
                in_dat_hld298[9:0] <= #DLY in_dat_wire298[9:0] ;
                in_dat_hld299[9:0] <= #DLY in_dat_wire299[9:0] ;
                in_dat_hld300[9:0] <= #DLY in_dat_wire300[9:0] ;
                in_dat_hld301[9:0] <= #DLY in_dat_wire301[9:0] ;
                in_dat_hld302[9:0] <= #DLY in_dat_wire302[9:0] ;
                in_dat_hld303[9:0] <= #DLY in_dat_wire303[9:0] ;
                in_dat_hld304[9:0] <= #DLY in_dat_wire304[9:0] ;
                in_dat_hld305[9:0] <= #DLY in_dat_wire305[9:0] ;
                in_dat_hld306[9:0] <= #DLY in_dat_wire306[9:0] ;
                in_dat_hld307[9:0] <= #DLY in_dat_wire307[9:0] ;
                in_dat_hld308[9:0] <= #DLY in_dat_wire308[9:0] ;
                in_dat_hld309[9:0] <= #DLY in_dat_wire309[9:0] ;
                in_dat_hld310[9:0] <= #DLY in_dat_wire310[9:0] ;
                in_dat_hld311[9:0] <= #DLY in_dat_wire311[9:0] ;
                in_dat_hld312[9:0] <= #DLY in_dat_wire312[9:0] ;
                in_dat_hld313[9:0] <= #DLY in_dat_wire313[9:0] ;
                in_dat_hld314[9:0] <= #DLY in_dat_wire314[9:0] ;
                in_dat_hld315[9:0] <= #DLY in_dat_wire315[9:0] ;
                in_dat_hld316[9:0] <= #DLY in_dat_wire316[9:0] ;
                in_dat_hld317[9:0] <= #DLY in_dat_wire317[9:0] ;
                in_dat_hld318[9:0] <= #DLY in_dat_wire318[9:0] ;
                in_dat_hld319[9:0] <= #DLY in_dat_wire319[9:0] ;
                in_dat_hld320[9:0] <= #DLY in_dat_wire320[9:0] ;
                in_dat_hld321[9:0] <= #DLY in_dat_wire321[9:0] ;
                in_dat_hld322[9:0] <= #DLY in_dat_wire322[9:0] ;
                in_dat_hld323[9:0] <= #DLY in_dat_wire323[9:0] ;
                in_dat_hld324[9:0] <= #DLY in_dat_wire324[9:0] ;
                in_dat_hld325[9:0] <= #DLY in_dat_wire325[9:0] ;
                in_dat_hld326[9:0] <= #DLY in_dat_wire326[9:0] ;
                in_dat_hld327[9:0] <= #DLY in_dat_wire327[9:0] ;
                in_dat_hld328[9:0] <= #DLY in_dat_wire328[9:0] ;
                in_dat_hld329[9:0] <= #DLY in_dat_wire329[9:0] ;
                in_dat_hld330[9:0] <= #DLY in_dat_wire330[9:0] ;
                in_dat_hld331[9:0] <= #DLY in_dat_wire331[9:0] ;
                in_dat_hld332[9:0] <= #DLY in_dat_wire332[9:0] ;
                in_dat_hld333[9:0] <= #DLY in_dat_wire333[9:0] ;
                in_dat_hld334[9:0] <= #DLY in_dat_wire334[9:0] ;
                in_dat_hld335[9:0] <= #DLY in_dat_wire335[9:0] ;
                in_dat_hld336[9:0] <= #DLY in_dat_wire336[9:0] ;
                in_dat_hld337[9:0] <= #DLY in_dat_wire337[9:0] ;
                in_dat_hld338[9:0] <= #DLY in_dat_wire338[9:0] ;
                in_dat_hld339[9:0] <= #DLY in_dat_wire339[9:0] ;
                in_dat_hld340[9:0] <= #DLY in_dat_wire340[9:0] ;
                in_dat_hld341[9:0] <= #DLY in_dat_wire341[9:0] ;
                in_dat_hld342[9:0] <= #DLY in_dat_wire342[9:0] ;
                in_dat_hld343[9:0] <= #DLY in_dat_wire343[9:0] ;
                in_dat_hld344[9:0] <= #DLY in_dat_wire344[9:0] ;
                in_dat_hld345[9:0] <= #DLY in_dat_wire345[9:0] ;
                in_dat_hld346[9:0] <= #DLY in_dat_wire346[9:0] ;
                in_dat_hld347[9:0] <= #DLY in_dat_wire347[9:0] ;
                in_dat_hld348[9:0] <= #DLY in_dat_wire348[9:0] ;
                in_dat_hld349[9:0] <= #DLY in_dat_wire349[9:0] ;
                in_dat_hld350[9:0] <= #DLY in_dat_wire350[9:0] ;
                in_dat_hld351[9:0] <= #DLY in_dat_wire351[9:0] ;
                in_dat_hld352[9:0] <= #DLY in_dat_wire352[9:0] ;
                in_dat_hld353[9:0] <= #DLY in_dat_wire353[9:0] ;
                in_dat_hld354[9:0] <= #DLY in_dat_wire354[9:0] ;
                in_dat_hld355[9:0] <= #DLY in_dat_wire355[9:0] ;
                in_dat_hld356[9:0] <= #DLY in_dat_wire356[9:0] ;
                in_dat_hld357[9:0] <= #DLY in_dat_wire357[9:0] ;
                in_dat_hld358[9:0] <= #DLY in_dat_wire358[9:0] ;
                in_dat_hld359[9:0] <= #DLY in_dat_wire359[9:0] ;
                in_dat_hld360[9:0] <= #DLY in_dat_wire360[9:0] ;
                in_dat_hld361[9:0] <= #DLY in_dat_wire361[9:0] ;
                in_dat_hld362[9:0] <= #DLY in_dat_wire362[9:0] ;
                in_dat_hld363[9:0] <= #DLY in_dat_wire363[9:0] ;
                in_dat_hld364[9:0] <= #DLY in_dat_wire364[9:0] ;
                in_dat_hld365[9:0] <= #DLY in_dat_wire365[9:0] ;
                in_dat_hld366[9:0] <= #DLY in_dat_wire366[9:0] ;
                in_dat_hld367[9:0] <= #DLY in_dat_wire367[9:0] ;
                in_dat_hld368[9:0] <= #DLY in_dat_wire368[9:0] ;
                in_dat_hld369[9:0] <= #DLY in_dat_wire369[9:0] ;
                in_dat_hld370[9:0] <= #DLY in_dat_wire370[9:0] ;
                in_dat_hld371[9:0] <= #DLY in_dat_wire371[9:0] ;
                in_dat_hld372[9:0] <= #DLY in_dat_wire372[9:0] ;
                in_dat_hld373[9:0] <= #DLY in_dat_wire373[9:0] ;
                in_dat_hld374[9:0] <= #DLY in_dat_wire374[9:0] ;
                in_dat_hld375[9:0] <= #DLY in_dat_wire375[9:0] ;
                in_dat_hld376[9:0] <= #DLY in_dat_wire376[9:0] ;
                in_dat_hld377[9:0] <= #DLY in_dat_wire377[9:0] ;
                in_dat_hld378[9:0] <= #DLY in_dat_wire378[9:0] ;
                in_dat_hld379[9:0] <= #DLY in_dat_wire379[9:0] ;
                in_dat_hld380[9:0] <= #DLY in_dat_wire380[9:0] ;
                in_dat_hld381[9:0] <= #DLY in_dat_wire381[9:0] ;
                in_dat_hld382[9:0] <= #DLY in_dat_wire382[9:0] ;
                in_dat_hld383[9:0] <= #DLY in_dat_wire383[9:0] ;
                in_dat_hld384[9:0] <= #DLY in_dat_wire384[9:0] ;
                in_dat_hld385[9:0] <= #DLY in_dat_wire385[9:0] ;
                in_dat_hld386[9:0] <= #DLY in_dat_wire386[9:0] ;
                in_dat_hld387[9:0] <= #DLY in_dat_wire387[9:0] ;
                in_dat_hld388[9:0] <= #DLY in_dat_wire388[9:0] ;
                in_dat_hld389[9:0] <= #DLY in_dat_wire389[9:0] ;
                in_dat_hld390[9:0] <= #DLY in_dat_wire390[9:0] ;
                in_dat_hld391[9:0] <= #DLY in_dat_wire391[9:0] ;
                in_dat_hld392[9:0] <= #DLY in_dat_wire392[9:0] ;
                in_dat_hld393[9:0] <= #DLY in_dat_wire393[9:0] ;
                in_dat_hld394[9:0] <= #DLY in_dat_wire394[9:0] ;
                in_dat_hld395[9:0] <= #DLY in_dat_wire395[9:0] ;
                in_dat_hld396[9:0] <= #DLY in_dat_wire396[9:0] ;
                in_dat_hld397[9:0] <= #DLY in_dat_wire397[9:0] ;
                in_dat_hld398[9:0] <= #DLY in_dat_wire398[9:0] ;
                in_dat_hld399[9:0] <= #DLY in_dat_wire399[9:0] ;
                in_dat_hld400[9:0] <= #DLY in_dat_wire400[9:0] ;
                in_dat_hld401[9:0] <= #DLY in_dat_wire401[9:0] ;
                in_dat_hld402[9:0] <= #DLY in_dat_wire402[9:0] ;
                in_dat_hld403[9:0] <= #DLY in_dat_wire403[9:0] ;
                in_dat_hld404[9:0] <= #DLY in_dat_wire404[9:0] ;
                in_dat_hld405[9:0] <= #DLY in_dat_wire405[9:0] ;
                in_dat_hld406[9:0] <= #DLY in_dat_wire406[9:0] ;
                in_dat_hld407[9:0] <= #DLY in_dat_wire407[9:0] ;
                in_dat_hld408[9:0] <= #DLY in_dat_wire408[9:0] ;
                in_dat_hld409[9:0] <= #DLY in_dat_wire409[9:0] ;
                in_dat_hld410[9:0] <= #DLY in_dat_wire410[9:0] ;
                in_dat_hld411[9:0] <= #DLY in_dat_wire411[9:0] ;
                in_dat_hld412[9:0] <= #DLY in_dat_wire412[9:0] ;
                in_dat_hld413[9:0] <= #DLY in_dat_wire413[9:0] ;
                in_dat_hld414[9:0] <= #DLY in_dat_wire414[9:0] ;
                in_dat_hld415[9:0] <= #DLY in_dat_wire415[9:0] ;
                in_dat_hld416[9:0] <= #DLY in_dat_wire416[9:0] ;
                in_dat_hld417[9:0] <= #DLY in_dat_wire417[9:0] ;
                in_dat_hld418[9:0] <= #DLY in_dat_wire418[9:0] ;
                in_dat_hld419[9:0] <= #DLY in_dat_wire419[9:0] ;
                in_dat_hld420[9:0] <= #DLY in_dat_wire420[9:0] ;
                in_dat_hld421[9:0] <= #DLY in_dat_wire421[9:0] ;
                in_dat_hld422[9:0] <= #DLY in_dat_wire422[9:0] ;
                in_dat_hld423[9:0] <= #DLY in_dat_wire423[9:0] ;
                in_dat_hld424[9:0] <= #DLY in_dat_wire424[9:0] ;
                in_dat_hld425[9:0] <= #DLY in_dat_wire425[9:0] ;
                in_dat_hld426[9:0] <= #DLY in_dat_wire426[9:0] ;
                in_dat_hld427[9:0] <= #DLY in_dat_wire427[9:0] ;
                in_dat_hld428[9:0] <= #DLY in_dat_wire428[9:0] ;
                in_dat_hld429[9:0] <= #DLY in_dat_wire429[9:0] ;
                in_dat_hld430[9:0] <= #DLY in_dat_wire430[9:0] ;
                in_dat_hld431[9:0] <= #DLY in_dat_wire431[9:0] ;
                in_dat_hld432[9:0] <= #DLY in_dat_wire432[9:0] ;
                in_dat_hld433[9:0] <= #DLY in_dat_wire433[9:0] ;
                in_dat_hld434[9:0] <= #DLY in_dat_wire434[9:0] ;
                in_dat_hld435[9:0] <= #DLY in_dat_wire435[9:0] ;
                in_dat_hld436[9:0] <= #DLY in_dat_wire436[9:0] ;
                in_dat_hld437[9:0] <= #DLY in_dat_wire437[9:0] ;
                in_dat_hld438[9:0] <= #DLY in_dat_wire438[9:0] ;
                in_dat_hld439[9:0] <= #DLY in_dat_wire439[9:0] ;
                in_dat_hld440[9:0] <= #DLY in_dat_wire440[9:0] ;
                in_dat_hld441[9:0] <= #DLY in_dat_wire441[9:0] ;
                in_dat_hld442[9:0] <= #DLY in_dat_wire442[9:0] ;
                in_dat_hld443[9:0] <= #DLY in_dat_wire443[9:0] ;
                in_dat_hld444[9:0] <= #DLY in_dat_wire444[9:0] ;
                in_dat_hld445[9:0] <= #DLY in_dat_wire445[9:0] ;
                in_dat_hld446[9:0] <= #DLY in_dat_wire446[9:0] ;
                in_dat_hld447[9:0] <= #DLY in_dat_wire447[9:0] ;
                in_dat_hld448[9:0] <= #DLY in_dat_wire448[9:0] ;
                in_dat_hld449[9:0] <= #DLY in_dat_wire449[9:0] ;
                in_dat_hld450[9:0] <= #DLY in_dat_wire450[9:0] ;
                in_dat_hld451[9:0] <= #DLY in_dat_wire451[9:0] ;
                in_dat_hld452[9:0] <= #DLY in_dat_wire452[9:0] ;
                in_dat_hld453[9:0] <= #DLY in_dat_wire453[9:0] ;
                in_dat_hld454[9:0] <= #DLY in_dat_wire454[9:0] ;
                in_dat_hld455[9:0] <= #DLY in_dat_wire455[9:0] ;
                in_dat_hld456[9:0] <= #DLY in_dat_wire456[9:0] ;
                in_dat_hld457[9:0] <= #DLY in_dat_wire457[9:0] ;
                in_dat_hld458[9:0] <= #DLY in_dat_wire458[9:0] ;
                in_dat_hld459[9:0] <= #DLY in_dat_wire459[9:0] ;
                in_dat_hld460[9:0] <= #DLY in_dat_wire460[9:0] ;
                in_dat_hld461[9:0] <= #DLY in_dat_wire461[9:0] ;
                in_dat_hld462[9:0] <= #DLY in_dat_wire462[9:0] ;
                in_dat_hld463[9:0] <= #DLY in_dat_wire463[9:0] ;
                in_dat_hld464[9:0] <= #DLY in_dat_wire464[9:0] ;
                in_dat_hld465[9:0] <= #DLY in_dat_wire465[9:0] ;
                in_dat_hld466[9:0] <= #DLY in_dat_wire466[9:0] ;
                in_dat_hld467[9:0] <= #DLY in_dat_wire467[9:0] ;
                in_dat_hld468[9:0] <= #DLY in_dat_wire468[9:0] ;
                in_dat_hld469[9:0] <= #DLY in_dat_wire469[9:0] ;
                in_dat_hld470[9:0] <= #DLY in_dat_wire470[9:0] ;
                in_dat_hld471[9:0] <= #DLY in_dat_wire471[9:0] ;
                in_dat_hld472[9:0] <= #DLY in_dat_wire472[9:0] ;
                in_dat_hld473[9:0] <= #DLY in_dat_wire473[9:0] ;
                in_dat_hld474[9:0] <= #DLY in_dat_wire474[9:0] ;
                in_dat_hld475[9:0] <= #DLY in_dat_wire475[9:0] ;
                in_dat_hld476[9:0] <= #DLY in_dat_wire476[9:0] ;
                in_dat_hld477[9:0] <= #DLY in_dat_wire477[9:0] ;
                in_dat_hld478[9:0] <= #DLY in_dat_wire478[9:0] ;
                in_dat_hld479[9:0] <= #DLY in_dat_wire479[9:0] ;
                in_dat_hld480[9:0] <= #DLY in_dat_wire480[9:0] ;
                in_dat_hld481[9:0] <= #DLY in_dat_wire481[9:0] ;
                in_dat_hld482[9:0] <= #DLY in_dat_wire482[9:0] ;
                in_dat_hld483[9:0] <= #DLY in_dat_wire483[9:0] ;
                in_dat_hld484[9:0] <= #DLY in_dat_wire484[9:0] ;
                in_dat_hld485[9:0] <= #DLY in_dat_wire485[9:0] ;
                in_dat_hld486[9:0] <= #DLY in_dat_wire486[9:0] ;
                in_dat_hld487[9:0] <= #DLY in_dat_wire487[9:0] ;
                in_dat_hld488[9:0] <= #DLY in_dat_wire488[9:0] ;
                in_dat_hld489[9:0] <= #DLY in_dat_wire489[9:0] ;
                in_dat_hld490[9:0] <= #DLY in_dat_wire490[9:0] ;
                in_dat_hld491[9:0] <= #DLY in_dat_wire491[9:0] ;
                in_dat_hld492[9:0] <= #DLY in_dat_wire492[9:0] ;
                in_dat_hld493[9:0] <= #DLY in_dat_wire493[9:0] ;
                in_dat_hld494[9:0] <= #DLY in_dat_wire494[9:0] ;
                in_dat_hld495[9:0] <= #DLY in_dat_wire495[9:0] ;
                in_dat_hld496[9:0] <= #DLY in_dat_wire496[9:0] ;
                in_dat_hld497[9:0] <= #DLY in_dat_wire497[9:0] ;
                in_dat_hld498[9:0] <= #DLY in_dat_wire498[9:0] ;
                in_dat_hld499[9:0] <= #DLY in_dat_wire499[9:0] ;
                in_dat_hld500[9:0] <= #DLY in_dat_wire500[9:0] ;
                in_dat_hld501[9:0] <= #DLY in_dat_wire501[9:0] ;
                in_dat_hld502[9:0] <= #DLY in_dat_wire502[9:0] ;
                in_dat_hld503[9:0] <= #DLY in_dat_wire503[9:0] ;
                in_dat_hld504[9:0] <= #DLY in_dat_wire504[9:0] ;
                in_dat_hld505[9:0] <= #DLY in_dat_wire505[9:0] ;
                in_dat_hld506[9:0] <= #DLY in_dat_wire506[9:0] ;
                in_dat_hld507[9:0] <= #DLY in_dat_wire507[9:0] ;
                in_dat_hld508[9:0] <= #DLY in_dat_wire508[9:0] ;
                in_dat_hld509[9:0] <= #DLY in_dat_wire509[9:0] ;
                in_dat_hld510[9:0] <= #DLY in_dat_wire510[9:0] ;
                in_dat_hld511[9:0] <= #DLY in_dat_wire511[9:0] ;
                in_dat_hld512[9:0] <= #DLY in_dat_wire512[9:0] ;
			end
		end
	end

    /****************************
    // pipeline[33] Active
    ****************************/
    wire [19:0] mult_wire01  = coe_dat_wire01[9:0]  * in_dat_hld01[9:0] ;
    wire [19:0] mult_wire02  = coe_dat_wire02[9:0]  * in_dat_hld02[9:0] ;
    wire [19:0] mult_wire03  = coe_dat_wire03[9:0]  * in_dat_hld03[9:0] ;
    wire [19:0] mult_wire04  = coe_dat_wire04[9:0]  * in_dat_hld04[9:0] ;
    wire [19:0] mult_wire05  = coe_dat_wire05[9:0]  * in_dat_hld05[9:0] ;
    wire [19:0] mult_wire06  = coe_dat_wire06[9:0]  * in_dat_hld06[9:0] ;
    wire [19:0] mult_wire07  = coe_dat_wire07[9:0]  * in_dat_hld07[9:0] ;
    wire [19:0] mult_wire08  = coe_dat_wire08[9:0]  * in_dat_hld08[9:0] ;
    wire [19:0] mult_wire09  = coe_dat_wire09[9:0]  * in_dat_hld09[9:0] ;
    wire [19:0] mult_wire10  = coe_dat_wire10[9:0]  * in_dat_hld10[9:0] ;
    wire [19:0] mult_wire11  = coe_dat_wire11[9:0]  * in_dat_hld11[9:0] ;
    wire [19:0] mult_wire12  = coe_dat_wire12[9:0]  * in_dat_hld12[9:0] ;
    wire [19:0] mult_wire13  = coe_dat_wire13[9:0]  * in_dat_hld13[9:0] ;
    wire [19:0] mult_wire14  = coe_dat_wire14[9:0]  * in_dat_hld14[9:0] ;
    wire [19:0] mult_wire15  = coe_dat_wire15[9:0]  * in_dat_hld15[9:0] ;
    wire [19:0] mult_wire16  = coe_dat_wire16[9:0]  * in_dat_hld16[9:0] ;
    wire [19:0] mult_wire17  = coe_dat_wire17[9:0]  * in_dat_hld17[9:0] ;
    wire [19:0] mult_wire18  = coe_dat_wire18[9:0]  * in_dat_hld18[9:0] ;
    wire [19:0] mult_wire19  = coe_dat_wire19[9:0]  * in_dat_hld19[9:0] ;
    wire [19:0] mult_wire20  = coe_dat_wire20[9:0]  * in_dat_hld20[9:0] ;
    wire [19:0] mult_wire21  = coe_dat_wire21[9:0]  * in_dat_hld21[9:0] ;
    wire [19:0] mult_wire22  = coe_dat_wire22[9:0]  * in_dat_hld22[9:0] ;
    wire [19:0] mult_wire23  = coe_dat_wire23[9:0]  * in_dat_hld23[9:0] ;
    wire [19:0] mult_wire24  = coe_dat_wire24[9:0]  * in_dat_hld24[9:0] ;
    wire [19:0] mult_wire25  = coe_dat_wire25[9:0]  * in_dat_hld25[9:0] ;
    wire [19:0] mult_wire26  = coe_dat_wire26[9:0]  * in_dat_hld26[9:0] ;
    wire [19:0] mult_wire27  = coe_dat_wire27[9:0]  * in_dat_hld27[9:0] ;
    wire [19:0] mult_wire28  = coe_dat_wire28[9:0]  * in_dat_hld28[9:0] ;
    wire [19:0] mult_wire29  = coe_dat_wire29[9:0]  * in_dat_hld29[9:0] ;
    wire [19:0] mult_wire30  = coe_dat_wire30[9:0]  * in_dat_hld30[9:0] ;
    wire [19:0] mult_wire31  = coe_dat_wire31[9:0]  * in_dat_hld31[9:0] ;
    wire [19:0] mult_wire32  = coe_dat_wire32[9:0]  * in_dat_hld32[9:0] ;
    wire [19:0] mult_wire33  = coe_dat_wire33[9:0]  * in_dat_hld33[9:0] ;
    wire [19:0] mult_wire34  = coe_dat_wire34[9:0]  * in_dat_hld34[9:0] ;
    wire [19:0] mult_wire35  = coe_dat_wire35[9:0]  * in_dat_hld35[9:0] ;
    wire [19:0] mult_wire36  = coe_dat_wire36[9:0]  * in_dat_hld36[9:0] ;
    wire [19:0] mult_wire37  = coe_dat_wire37[9:0]  * in_dat_hld37[9:0] ;
    wire [19:0] mult_wire38  = coe_dat_wire38[9:0]  * in_dat_hld38[9:0] ;
    wire [19:0] mult_wire39  = coe_dat_wire39[9:0]  * in_dat_hld39[9:0] ;
    wire [19:0] mult_wire40  = coe_dat_wire40[9:0]  * in_dat_hld40[9:0] ;
    wire [19:0] mult_wire41  = coe_dat_wire41[9:0]  * in_dat_hld41[9:0] ;
    wire [19:0] mult_wire42  = coe_dat_wire42[9:0]  * in_dat_hld42[9:0] ;
    wire [19:0] mult_wire43  = coe_dat_wire43[9:0]  * in_dat_hld43[9:0] ;
    wire [19:0] mult_wire44  = coe_dat_wire44[9:0]  * in_dat_hld44[9:0] ;
    wire [19:0] mult_wire45  = coe_dat_wire45[9:0]  * in_dat_hld45[9:0] ;
    wire [19:0] mult_wire46  = coe_dat_wire46[9:0]  * in_dat_hld46[9:0] ;
    wire [19:0] mult_wire47  = coe_dat_wire47[9:0]  * in_dat_hld47[9:0] ;
    wire [19:0] mult_wire48  = coe_dat_wire48[9:0]  * in_dat_hld48[9:0] ;
    wire [19:0] mult_wire49  = coe_dat_wire49[9:0]  * in_dat_hld49[9:0] ;
    wire [19:0] mult_wire50  = coe_dat_wire50[9:0]  * in_dat_hld50[9:0] ;
    wire [19:0] mult_wire51  = coe_dat_wire51[9:0]  * in_dat_hld51[9:0] ;
    wire [19:0] mult_wire52  = coe_dat_wire52[9:0]  * in_dat_hld52[9:0] ;
    wire [19:0] mult_wire53  = coe_dat_wire53[9:0]  * in_dat_hld53[9:0] ;
    wire [19:0] mult_wire54  = coe_dat_wire54[9:0]  * in_dat_hld54[9:0] ;
    wire [19:0] mult_wire55  = coe_dat_wire55[9:0]  * in_dat_hld55[9:0] ;
    wire [19:0] mult_wire56  = coe_dat_wire56[9:0]  * in_dat_hld56[9:0] ;
    wire [19:0] mult_wire57  = coe_dat_wire57[9:0]  * in_dat_hld57[9:0] ;
    wire [19:0] mult_wire58  = coe_dat_wire58[9:0]  * in_dat_hld58[9:0] ;
    wire [19:0] mult_wire59  = coe_dat_wire59[9:0]  * in_dat_hld59[9:0] ;
    wire [19:0] mult_wire60  = coe_dat_wire60[9:0]  * in_dat_hld60[9:0] ;
    wire [19:0] mult_wire61  = coe_dat_wire61[9:0]  * in_dat_hld61[9:0] ;
    wire [19:0] mult_wire62  = coe_dat_wire62[9:0]  * in_dat_hld62[9:0] ;
    wire [19:0] mult_wire63  = coe_dat_wire63[9:0]  * in_dat_hld63[9:0] ;
    wire [19:0] mult_wire64  = coe_dat_wire64[9:0]  * in_dat_hld64[9:0] ;
    wire [19:0] mult_wire65  = coe_dat_wire65[9:0]  * in_dat_hld65[9:0] ;
    wire [19:0] mult_wire66  = coe_dat_wire66[9:0]  * in_dat_hld66[9:0] ;
    wire [19:0] mult_wire67  = coe_dat_wire67[9:0]  * in_dat_hld67[9:0] ;
    wire [19:0] mult_wire68  = coe_dat_wire68[9:0]  * in_dat_hld68[9:0] ;
    wire [19:0] mult_wire69  = coe_dat_wire69[9:0]  * in_dat_hld69[9:0] ;
    wire [19:0] mult_wire70  = coe_dat_wire70[9:0]  * in_dat_hld70[9:0] ;
    wire [19:0] mult_wire71  = coe_dat_wire71[9:0]  * in_dat_hld71[9:0] ;
    wire [19:0] mult_wire72  = coe_dat_wire72[9:0]  * in_dat_hld72[9:0] ;
    wire [19:0] mult_wire73  = coe_dat_wire73[9:0]  * in_dat_hld73[9:0] ;
    wire [19:0] mult_wire74  = coe_dat_wire74[9:0]  * in_dat_hld74[9:0] ;
    wire [19:0] mult_wire75  = coe_dat_wire75[9:0]  * in_dat_hld75[9:0] ;
    wire [19:0] mult_wire76  = coe_dat_wire76[9:0]  * in_dat_hld76[9:0] ;
    wire [19:0] mult_wire77  = coe_dat_wire77[9:0]  * in_dat_hld77[9:0] ;
    wire [19:0] mult_wire78  = coe_dat_wire78[9:0]  * in_dat_hld78[9:0] ;
    wire [19:0] mult_wire79  = coe_dat_wire79[9:0]  * in_dat_hld79[9:0] ;
    wire [19:0] mult_wire80  = coe_dat_wire80[9:0]  * in_dat_hld80[9:0] ;
    wire [19:0] mult_wire81  = coe_dat_wire81[9:0]  * in_dat_hld81[9:0] ;
    wire [19:0] mult_wire82  = coe_dat_wire82[9:0]  * in_dat_hld82[9:0] ;
    wire [19:0] mult_wire83  = coe_dat_wire83[9:0]  * in_dat_hld83[9:0] ;
    wire [19:0] mult_wire84  = coe_dat_wire84[9:0]  * in_dat_hld84[9:0] ;
    wire [19:0] mult_wire85  = coe_dat_wire85[9:0]  * in_dat_hld85[9:0] ;
    wire [19:0] mult_wire86  = coe_dat_wire86[9:0]  * in_dat_hld86[9:0] ;
    wire [19:0] mult_wire87  = coe_dat_wire87[9:0]  * in_dat_hld87[9:0] ;
    wire [19:0] mult_wire88  = coe_dat_wire88[9:0]  * in_dat_hld88[9:0] ;
    wire [19:0] mult_wire89  = coe_dat_wire89[9:0]  * in_dat_hld89[9:0] ;
    wire [19:0] mult_wire90  = coe_dat_wire90[9:0]  * in_dat_hld90[9:0] ;
    wire [19:0] mult_wire91  = coe_dat_wire91[9:0]  * in_dat_hld91[9:0] ;
    wire [19:0] mult_wire92  = coe_dat_wire92[9:0]  * in_dat_hld92[9:0] ;
    wire [19:0] mult_wire93  = coe_dat_wire93[9:0]  * in_dat_hld93[9:0] ;
    wire [19:0] mult_wire94  = coe_dat_wire94[9:0]  * in_dat_hld94[9:0] ;
    wire [19:0] mult_wire95  = coe_dat_wire95[9:0]  * in_dat_hld95[9:0] ;
    wire [19:0] mult_wire96  = coe_dat_wire96[9:0]  * in_dat_hld96[9:0] ;
    wire [19:0] mult_wire97  = coe_dat_wire97[9:0]  * in_dat_hld97[9:0] ;
    wire [19:0] mult_wire98  = coe_dat_wire98[9:0]  * in_dat_hld98[9:0] ;
    wire [19:0] mult_wire99  = coe_dat_wire99[9:0]  * in_dat_hld99[9:0] ;
    wire [19:0] mult_wire100 = coe_dat_wire100[9:0] * in_dat_hld100[9:0] ;
    wire [19:0] mult_wire101 = coe_dat_wire101[9:0] * in_dat_hld101[9:0] ;
    wire [19:0] mult_wire102 = coe_dat_wire102[9:0] * in_dat_hld102[9:0] ;
    wire [19:0] mult_wire103 = coe_dat_wire103[9:0] * in_dat_hld103[9:0] ;
    wire [19:0] mult_wire104 = coe_dat_wire104[9:0] * in_dat_hld104[9:0] ;
    wire [19:0] mult_wire105 = coe_dat_wire105[9:0] * in_dat_hld105[9:0] ;
    wire [19:0] mult_wire106 = coe_dat_wire106[9:0] * in_dat_hld106[9:0] ;
    wire [19:0] mult_wire107 = coe_dat_wire107[9:0] * in_dat_hld107[9:0] ;
    wire [19:0] mult_wire108 = coe_dat_wire108[9:0] * in_dat_hld108[9:0] ;
    wire [19:0] mult_wire109 = coe_dat_wire109[9:0] * in_dat_hld109[9:0] ;
    wire [19:0] mult_wire110 = coe_dat_wire110[9:0] * in_dat_hld110[9:0] ;
    wire [19:0] mult_wire111 = coe_dat_wire111[9:0] * in_dat_hld111[9:0] ;
    wire [19:0] mult_wire112 = coe_dat_wire112[9:0] * in_dat_hld112[9:0] ;
    wire [19:0] mult_wire113 = coe_dat_wire113[9:0] * in_dat_hld113[9:0] ;
    wire [19:0] mult_wire114 = coe_dat_wire114[9:0] * in_dat_hld114[9:0] ;
    wire [19:0] mult_wire115 = coe_dat_wire115[9:0] * in_dat_hld115[9:0] ;
    wire [19:0] mult_wire116 = coe_dat_wire116[9:0] * in_dat_hld116[9:0] ;
    wire [19:0] mult_wire117 = coe_dat_wire117[9:0] * in_dat_hld117[9:0] ;
    wire [19:0] mult_wire118 = coe_dat_wire118[9:0] * in_dat_hld118[9:0] ;
    wire [19:0] mult_wire119 = coe_dat_wire119[9:0] * in_dat_hld119[9:0] ;
    wire [19:0] mult_wire120 = coe_dat_wire120[9:0] * in_dat_hld120[9:0] ;
    wire [19:0] mult_wire121 = coe_dat_wire121[9:0] * in_dat_hld121[9:0] ;
    wire [19:0] mult_wire122 = coe_dat_wire122[9:0] * in_dat_hld122[9:0] ;
    wire [19:0] mult_wire123 = coe_dat_wire123[9:0] * in_dat_hld123[9:0] ;
    wire [19:0] mult_wire124 = coe_dat_wire124[9:0] * in_dat_hld124[9:0] ;
    wire [19:0] mult_wire125 = coe_dat_wire125[9:0] * in_dat_hld125[9:0] ;
    wire [19:0] mult_wire126 = coe_dat_wire126[9:0] * in_dat_hld126[9:0] ;
    wire [19:0] mult_wire127 = coe_dat_wire127[9:0] * in_dat_hld127[9:0] ;
    wire [19:0] mult_wire128 = coe_dat_wire128[9:0] * in_dat_hld128[9:0] ;
    wire [19:0] mult_wire129 = coe_dat_wire129[9:0] * in_dat_hld129[9:0] ;
    wire [19:0] mult_wire130 = coe_dat_wire130[9:0] * in_dat_hld130[9:0] ;
    wire [19:0] mult_wire131 = coe_dat_wire131[9:0] * in_dat_hld131[9:0] ;
    wire [19:0] mult_wire132 = coe_dat_wire132[9:0] * in_dat_hld132[9:0] ;
    wire [19:0] mult_wire133 = coe_dat_wire133[9:0] * in_dat_hld133[9:0] ;
    wire [19:0] mult_wire134 = coe_dat_wire134[9:0] * in_dat_hld134[9:0] ;
    wire [19:0] mult_wire135 = coe_dat_wire135[9:0] * in_dat_hld135[9:0] ;
    wire [19:0] mult_wire136 = coe_dat_wire136[9:0] * in_dat_hld136[9:0] ;
    wire [19:0] mult_wire137 = coe_dat_wire137[9:0] * in_dat_hld137[9:0] ;
    wire [19:0] mult_wire138 = coe_dat_wire138[9:0] * in_dat_hld138[9:0] ;
    wire [19:0] mult_wire139 = coe_dat_wire139[9:0] * in_dat_hld139[9:0] ;
    wire [19:0] mult_wire140 = coe_dat_wire140[9:0] * in_dat_hld140[9:0] ;
    wire [19:0] mult_wire141 = coe_dat_wire141[9:0] * in_dat_hld141[9:0] ;
    wire [19:0] mult_wire142 = coe_dat_wire142[9:0] * in_dat_hld142[9:0] ;
    wire [19:0] mult_wire143 = coe_dat_wire143[9:0] * in_dat_hld143[9:0] ;
    wire [19:0] mult_wire144 = coe_dat_wire144[9:0] * in_dat_hld144[9:0] ;
    wire [19:0] mult_wire145 = coe_dat_wire145[9:0] * in_dat_hld145[9:0] ;
    wire [19:0] mult_wire146 = coe_dat_wire146[9:0] * in_dat_hld146[9:0] ;
    wire [19:0] mult_wire147 = coe_dat_wire147[9:0] * in_dat_hld147[9:0] ;
    wire [19:0] mult_wire148 = coe_dat_wire148[9:0] * in_dat_hld148[9:0] ;
    wire [19:0] mult_wire149 = coe_dat_wire149[9:0] * in_dat_hld149[9:0] ;
    wire [19:0] mult_wire150 = coe_dat_wire150[9:0] * in_dat_hld150[9:0] ;
    wire [19:0] mult_wire151 = coe_dat_wire151[9:0] * in_dat_hld151[9:0] ;
    wire [19:0] mult_wire152 = coe_dat_wire152[9:0] * in_dat_hld152[9:0] ;
    wire [19:0] mult_wire153 = coe_dat_wire153[9:0] * in_dat_hld153[9:0] ;
    wire [19:0] mult_wire154 = coe_dat_wire154[9:0] * in_dat_hld154[9:0] ;
    wire [19:0] mult_wire155 = coe_dat_wire155[9:0] * in_dat_hld155[9:0] ;
    wire [19:0] mult_wire156 = coe_dat_wire156[9:0] * in_dat_hld156[9:0] ;
    wire [19:0] mult_wire157 = coe_dat_wire157[9:0] * in_dat_hld157[9:0] ;
    wire [19:0] mult_wire158 = coe_dat_wire158[9:0] * in_dat_hld158[9:0] ;
    wire [19:0] mult_wire159 = coe_dat_wire159[9:0] * in_dat_hld159[9:0] ;
    wire [19:0] mult_wire160 = coe_dat_wire160[9:0] * in_dat_hld160[9:0] ;
    wire [19:0] mult_wire161 = coe_dat_wire161[9:0] * in_dat_hld161[9:0] ;
    wire [19:0] mult_wire162 = coe_dat_wire162[9:0] * in_dat_hld162[9:0] ;
    wire [19:0] mult_wire163 = coe_dat_wire163[9:0] * in_dat_hld163[9:0] ;
    wire [19:0] mult_wire164 = coe_dat_wire164[9:0] * in_dat_hld164[9:0] ;
    wire [19:0] mult_wire165 = coe_dat_wire165[9:0] * in_dat_hld165[9:0] ;
    wire [19:0] mult_wire166 = coe_dat_wire166[9:0] * in_dat_hld166[9:0] ;
    wire [19:0] mult_wire167 = coe_dat_wire167[9:0] * in_dat_hld167[9:0] ;
    wire [19:0] mult_wire168 = coe_dat_wire168[9:0] * in_dat_hld168[9:0] ;
    wire [19:0] mult_wire169 = coe_dat_wire169[9:0] * in_dat_hld169[9:0] ;
    wire [19:0] mult_wire170 = coe_dat_wire170[9:0] * in_dat_hld170[9:0] ;
    wire [19:0] mult_wire171 = coe_dat_wire171[9:0] * in_dat_hld171[9:0] ;
    wire [19:0] mult_wire172 = coe_dat_wire172[9:0] * in_dat_hld172[9:0] ;
    wire [19:0] mult_wire173 = coe_dat_wire173[9:0] * in_dat_hld173[9:0] ;
    wire [19:0] mult_wire174 = coe_dat_wire174[9:0] * in_dat_hld174[9:0] ;
    wire [19:0] mult_wire175 = coe_dat_wire175[9:0] * in_dat_hld175[9:0] ;
    wire [19:0] mult_wire176 = coe_dat_wire176[9:0] * in_dat_hld176[9:0] ;
    wire [19:0] mult_wire177 = coe_dat_wire177[9:0] * in_dat_hld177[9:0] ;
    wire [19:0] mult_wire178 = coe_dat_wire178[9:0] * in_dat_hld178[9:0] ;
    wire [19:0] mult_wire179 = coe_dat_wire179[9:0] * in_dat_hld179[9:0] ;
    wire [19:0] mult_wire180 = coe_dat_wire180[9:0] * in_dat_hld180[9:0] ;
    wire [19:0] mult_wire181 = coe_dat_wire181[9:0] * in_dat_hld181[9:0] ;
    wire [19:0] mult_wire182 = coe_dat_wire182[9:0] * in_dat_hld182[9:0] ;
    wire [19:0] mult_wire183 = coe_dat_wire183[9:0] * in_dat_hld183[9:0] ;
    wire [19:0] mult_wire184 = coe_dat_wire184[9:0] * in_dat_hld184[9:0] ;
    wire [19:0] mult_wire185 = coe_dat_wire185[9:0] * in_dat_hld185[9:0] ;
    wire [19:0] mult_wire186 = coe_dat_wire186[9:0] * in_dat_hld186[9:0] ;
    wire [19:0] mult_wire187 = coe_dat_wire187[9:0] * in_dat_hld187[9:0] ;
    wire [19:0] mult_wire188 = coe_dat_wire188[9:0] * in_dat_hld188[9:0] ;
    wire [19:0] mult_wire189 = coe_dat_wire189[9:0] * in_dat_hld189[9:0] ;
    wire [19:0] mult_wire190 = coe_dat_wire190[9:0] * in_dat_hld190[9:0] ;
    wire [19:0] mult_wire191 = coe_dat_wire191[9:0] * in_dat_hld191[9:0] ;
    wire [19:0] mult_wire192 = coe_dat_wire192[9:0] * in_dat_hld192[9:0] ;
    wire [19:0] mult_wire193 = coe_dat_wire193[9:0] * in_dat_hld193[9:0] ;
    wire [19:0] mult_wire194 = coe_dat_wire194[9:0] * in_dat_hld194[9:0] ;
    wire [19:0] mult_wire195 = coe_dat_wire195[9:0] * in_dat_hld195[9:0] ;
    wire [19:0] mult_wire196 = coe_dat_wire196[9:0] * in_dat_hld196[9:0] ;
    wire [19:0] mult_wire197 = coe_dat_wire197[9:0] * in_dat_hld197[9:0] ;
    wire [19:0] mult_wire198 = coe_dat_wire198[9:0] * in_dat_hld198[9:0] ;
    wire [19:0] mult_wire199 = coe_dat_wire199[9:0] * in_dat_hld199[9:0] ;
    wire [19:0] mult_wire200 = coe_dat_wire200[9:0] * in_dat_hld200[9:0] ;
    wire [19:0] mult_wire201 = coe_dat_wire201[9:0] * in_dat_hld201[9:0] ;
    wire [19:0] mult_wire202 = coe_dat_wire202[9:0] * in_dat_hld202[9:0] ;
    wire [19:0] mult_wire203 = coe_dat_wire203[9:0] * in_dat_hld203[9:0] ;
    wire [19:0] mult_wire204 = coe_dat_wire204[9:0] * in_dat_hld204[9:0] ;
    wire [19:0] mult_wire205 = coe_dat_wire205[9:0] * in_dat_hld205[9:0] ;
    wire [19:0] mult_wire206 = coe_dat_wire206[9:0] * in_dat_hld206[9:0] ;
    wire [19:0] mult_wire207 = coe_dat_wire207[9:0] * in_dat_hld207[9:0] ;
    wire [19:0] mult_wire208 = coe_dat_wire208[9:0] * in_dat_hld208[9:0] ;
    wire [19:0] mult_wire209 = coe_dat_wire209[9:0] * in_dat_hld209[9:0] ;
    wire [19:0] mult_wire210 = coe_dat_wire210[9:0] * in_dat_hld210[9:0] ;
    wire [19:0] mult_wire211 = coe_dat_wire211[9:0] * in_dat_hld211[9:0] ;
    wire [19:0] mult_wire212 = coe_dat_wire212[9:0] * in_dat_hld212[9:0] ;
    wire [19:0] mult_wire213 = coe_dat_wire213[9:0] * in_dat_hld213[9:0] ;
    wire [19:0] mult_wire214 = coe_dat_wire214[9:0] * in_dat_hld214[9:0] ;
    wire [19:0] mult_wire215 = coe_dat_wire215[9:0] * in_dat_hld215[9:0] ;
    wire [19:0] mult_wire216 = coe_dat_wire216[9:0] * in_dat_hld216[9:0] ;
    wire [19:0] mult_wire217 = coe_dat_wire217[9:0] * in_dat_hld217[9:0] ;
    wire [19:0] mult_wire218 = coe_dat_wire218[9:0] * in_dat_hld218[9:0] ;
    wire [19:0] mult_wire219 = coe_dat_wire219[9:0] * in_dat_hld219[9:0] ;
    wire [19:0] mult_wire220 = coe_dat_wire220[9:0] * in_dat_hld220[9:0] ;
    wire [19:0] mult_wire221 = coe_dat_wire221[9:0] * in_dat_hld221[9:0] ;
    wire [19:0] mult_wire222 = coe_dat_wire222[9:0] * in_dat_hld222[9:0] ;
    wire [19:0] mult_wire223 = coe_dat_wire223[9:0] * in_dat_hld223[9:0] ;
    wire [19:0] mult_wire224 = coe_dat_wire224[9:0] * in_dat_hld224[9:0] ;
    wire [19:0] mult_wire225 = coe_dat_wire225[9:0] * in_dat_hld225[9:0] ;
    wire [19:0] mult_wire226 = coe_dat_wire226[9:0] * in_dat_hld226[9:0] ;
    wire [19:0] mult_wire227 = coe_dat_wire227[9:0] * in_dat_hld227[9:0] ;
    wire [19:0] mult_wire228 = coe_dat_wire228[9:0] * in_dat_hld228[9:0] ;
    wire [19:0] mult_wire229 = coe_dat_wire229[9:0] * in_dat_hld229[9:0] ;
    wire [19:0] mult_wire230 = coe_dat_wire230[9:0] * in_dat_hld230[9:0] ;
    wire [19:0] mult_wire231 = coe_dat_wire231[9:0] * in_dat_hld231[9:0] ;
    wire [19:0] mult_wire232 = coe_dat_wire232[9:0] * in_dat_hld232[9:0] ;
    wire [19:0] mult_wire233 = coe_dat_wire233[9:0] * in_dat_hld233[9:0] ;
    wire [19:0] mult_wire234 = coe_dat_wire234[9:0] * in_dat_hld234[9:0] ;
    wire [19:0] mult_wire235 = coe_dat_wire235[9:0] * in_dat_hld235[9:0] ;
    wire [19:0] mult_wire236 = coe_dat_wire236[9:0] * in_dat_hld236[9:0] ;
    wire [19:0] mult_wire237 = coe_dat_wire237[9:0] * in_dat_hld237[9:0] ;
    wire [19:0] mult_wire238 = coe_dat_wire238[9:0] * in_dat_hld238[9:0] ;
    wire [19:0] mult_wire239 = coe_dat_wire239[9:0] * in_dat_hld239[9:0] ;
    wire [19:0] mult_wire240 = coe_dat_wire240[9:0] * in_dat_hld240[9:0] ;
    wire [19:0] mult_wire241 = coe_dat_wire241[9:0] * in_dat_hld241[9:0] ;
    wire [19:0] mult_wire242 = coe_dat_wire242[9:0] * in_dat_hld242[9:0] ;
    wire [19:0] mult_wire243 = coe_dat_wire243[9:0] * in_dat_hld243[9:0] ;
    wire [19:0] mult_wire244 = coe_dat_wire244[9:0] * in_dat_hld244[9:0] ;
    wire [19:0] mult_wire245 = coe_dat_wire245[9:0] * in_dat_hld245[9:0] ;
    wire [19:0] mult_wire246 = coe_dat_wire246[9:0] * in_dat_hld246[9:0] ;
    wire [19:0] mult_wire247 = coe_dat_wire247[9:0] * in_dat_hld247[9:0] ;
    wire [19:0] mult_wire248 = coe_dat_wire248[9:0] * in_dat_hld248[9:0] ;
    wire [19:0] mult_wire249 = coe_dat_wire249[9:0] * in_dat_hld249[9:0] ;
    wire [19:0] mult_wire250 = coe_dat_wire250[9:0] * in_dat_hld250[9:0] ;
    wire [19:0] mult_wire251 = coe_dat_wire251[9:0] * in_dat_hld251[9:0] ;
    wire [19:0] mult_wire252 = coe_dat_wire252[9:0] * in_dat_hld252[9:0] ;
    wire [19:0] mult_wire253 = coe_dat_wire253[9:0] * in_dat_hld253[9:0] ;
    wire [19:0] mult_wire254 = coe_dat_wire254[9:0] * in_dat_hld254[9:0] ;
    wire [19:0] mult_wire255 = coe_dat_wire255[9:0] * in_dat_hld255[9:0] ;
    wire [19:0] mult_wire256 = coe_dat_wire256[9:0] * in_dat_hld256[9:0] ;
    wire [19:0] mult_wire257 = coe_dat_wire257[9:0] * in_dat_hld257[9:0] ;
    wire [19:0] mult_wire258 = coe_dat_wire258[9:0] * in_dat_hld258[9:0] ;
    wire [19:0] mult_wire259 = coe_dat_wire259[9:0] * in_dat_hld259[9:0] ;
    wire [19:0] mult_wire260 = coe_dat_wire260[9:0] * in_dat_hld260[9:0] ;
    wire [19:0] mult_wire261 = coe_dat_wire261[9:0] * in_dat_hld261[9:0] ;
    wire [19:0] mult_wire262 = coe_dat_wire262[9:0] * in_dat_hld262[9:0] ;
    wire [19:0] mult_wire263 = coe_dat_wire263[9:0] * in_dat_hld263[9:0] ;
    wire [19:0] mult_wire264 = coe_dat_wire264[9:0] * in_dat_hld264[9:0] ;
    wire [19:0] mult_wire265 = coe_dat_wire265[9:0] * in_dat_hld265[9:0] ;
    wire [19:0] mult_wire266 = coe_dat_wire266[9:0] * in_dat_hld266[9:0] ;
    wire [19:0] mult_wire267 = coe_dat_wire267[9:0] * in_dat_hld267[9:0] ;
    wire [19:0] mult_wire268 = coe_dat_wire268[9:0] * in_dat_hld268[9:0] ;
    wire [19:0] mult_wire269 = coe_dat_wire269[9:0] * in_dat_hld269[9:0] ;
    wire [19:0] mult_wire270 = coe_dat_wire270[9:0] * in_dat_hld270[9:0] ;
    wire [19:0] mult_wire271 = coe_dat_wire271[9:0] * in_dat_hld271[9:0] ;
    wire [19:0] mult_wire272 = coe_dat_wire272[9:0] * in_dat_hld272[9:0] ;
    wire [19:0] mult_wire273 = coe_dat_wire273[9:0] * in_dat_hld273[9:0] ;
    wire [19:0] mult_wire274 = coe_dat_wire274[9:0] * in_dat_hld274[9:0] ;
    wire [19:0] mult_wire275 = coe_dat_wire275[9:0] * in_dat_hld275[9:0] ;
    wire [19:0] mult_wire276 = coe_dat_wire276[9:0] * in_dat_hld276[9:0] ;
    wire [19:0] mult_wire277 = coe_dat_wire277[9:0] * in_dat_hld277[9:0] ;
    wire [19:0] mult_wire278 = coe_dat_wire278[9:0] * in_dat_hld278[9:0] ;
    wire [19:0] mult_wire279 = coe_dat_wire279[9:0] * in_dat_hld279[9:0] ;
    wire [19:0] mult_wire280 = coe_dat_wire280[9:0] * in_dat_hld280[9:0] ;
    wire [19:0] mult_wire281 = coe_dat_wire281[9:0] * in_dat_hld281[9:0] ;
    wire [19:0] mult_wire282 = coe_dat_wire282[9:0] * in_dat_hld282[9:0] ;
    wire [19:0] mult_wire283 = coe_dat_wire283[9:0] * in_dat_hld283[9:0] ;
    wire [19:0] mult_wire284 = coe_dat_wire284[9:0] * in_dat_hld284[9:0] ;
    wire [19:0] mult_wire285 = coe_dat_wire285[9:0] * in_dat_hld285[9:0] ;
    wire [19:0] mult_wire286 = coe_dat_wire286[9:0] * in_dat_hld286[9:0] ;
    wire [19:0] mult_wire287 = coe_dat_wire287[9:0] * in_dat_hld287[9:0] ;
    wire [19:0] mult_wire288 = coe_dat_wire288[9:0] * in_dat_hld288[9:0] ;
    wire [19:0] mult_wire289 = coe_dat_wire289[9:0] * in_dat_hld289[9:0] ;
    wire [19:0] mult_wire290 = coe_dat_wire290[9:0] * in_dat_hld290[9:0] ;
    wire [19:0] mult_wire291 = coe_dat_wire291[9:0] * in_dat_hld291[9:0] ;
    wire [19:0] mult_wire292 = coe_dat_wire292[9:0] * in_dat_hld292[9:0] ;
    wire [19:0] mult_wire293 = coe_dat_wire293[9:0] * in_dat_hld293[9:0] ;
    wire [19:0] mult_wire294 = coe_dat_wire294[9:0] * in_dat_hld294[9:0] ;
    wire [19:0] mult_wire295 = coe_dat_wire295[9:0] * in_dat_hld295[9:0] ;
    wire [19:0] mult_wire296 = coe_dat_wire296[9:0] * in_dat_hld296[9:0] ;
    wire [19:0] mult_wire297 = coe_dat_wire297[9:0] * in_dat_hld297[9:0] ;
    wire [19:0] mult_wire298 = coe_dat_wire298[9:0] * in_dat_hld298[9:0] ;
    wire [19:0] mult_wire299 = coe_dat_wire299[9:0] * in_dat_hld299[9:0] ;
    wire [19:0] mult_wire300 = coe_dat_wire300[9:0] * in_dat_hld300[9:0] ;
    wire [19:0] mult_wire301 = coe_dat_wire301[9:0] * in_dat_hld301[9:0] ;
    wire [19:0] mult_wire302 = coe_dat_wire302[9:0] * in_dat_hld302[9:0] ;
    wire [19:0] mult_wire303 = coe_dat_wire303[9:0] * in_dat_hld303[9:0] ;
    wire [19:0] mult_wire304 = coe_dat_wire304[9:0] * in_dat_hld304[9:0] ;
    wire [19:0] mult_wire305 = coe_dat_wire305[9:0] * in_dat_hld305[9:0] ;
    wire [19:0] mult_wire306 = coe_dat_wire306[9:0] * in_dat_hld306[9:0] ;
    wire [19:0] mult_wire307 = coe_dat_wire307[9:0] * in_dat_hld307[9:0] ;
    wire [19:0] mult_wire308 = coe_dat_wire308[9:0] * in_dat_hld308[9:0] ;
    wire [19:0] mult_wire309 = coe_dat_wire309[9:0] * in_dat_hld309[9:0] ;
    wire [19:0] mult_wire310 = coe_dat_wire310[9:0] * in_dat_hld310[9:0] ;
    wire [19:0] mult_wire311 = coe_dat_wire311[9:0] * in_dat_hld311[9:0] ;
    wire [19:0] mult_wire312 = coe_dat_wire312[9:0] * in_dat_hld312[9:0] ;
    wire [19:0] mult_wire313 = coe_dat_wire313[9:0] * in_dat_hld313[9:0] ;
    wire [19:0] mult_wire314 = coe_dat_wire314[9:0] * in_dat_hld314[9:0] ;
    wire [19:0] mult_wire315 = coe_dat_wire315[9:0] * in_dat_hld315[9:0] ;
    wire [19:0] mult_wire316 = coe_dat_wire316[9:0] * in_dat_hld316[9:0] ;
    wire [19:0] mult_wire317 = coe_dat_wire317[9:0] * in_dat_hld317[9:0] ;
    wire [19:0] mult_wire318 = coe_dat_wire318[9:0] * in_dat_hld318[9:0] ;
    wire [19:0] mult_wire319 = coe_dat_wire319[9:0] * in_dat_hld319[9:0] ;
    wire [19:0] mult_wire320 = coe_dat_wire320[9:0] * in_dat_hld320[9:0] ;
    wire [19:0] mult_wire321 = coe_dat_wire321[9:0] * in_dat_hld321[9:0] ;
    wire [19:0] mult_wire322 = coe_dat_wire322[9:0] * in_dat_hld322[9:0] ;
    wire [19:0] mult_wire323 = coe_dat_wire323[9:0] * in_dat_hld323[9:0] ;
    wire [19:0] mult_wire324 = coe_dat_wire324[9:0] * in_dat_hld324[9:0] ;
    wire [19:0] mult_wire325 = coe_dat_wire325[9:0] * in_dat_hld325[9:0] ;
    wire [19:0] mult_wire326 = coe_dat_wire326[9:0] * in_dat_hld326[9:0] ;
    wire [19:0] mult_wire327 = coe_dat_wire327[9:0] * in_dat_hld327[9:0] ;
    wire [19:0] mult_wire328 = coe_dat_wire328[9:0] * in_dat_hld328[9:0] ;
    wire [19:0] mult_wire329 = coe_dat_wire329[9:0] * in_dat_hld329[9:0] ;
    wire [19:0] mult_wire330 = coe_dat_wire330[9:0] * in_dat_hld330[9:0] ;
    wire [19:0] mult_wire331 = coe_dat_wire331[9:0] * in_dat_hld331[9:0] ;
    wire [19:0] mult_wire332 = coe_dat_wire332[9:0] * in_dat_hld332[9:0] ;
    wire [19:0] mult_wire333 = coe_dat_wire333[9:0] * in_dat_hld333[9:0] ;
    wire [19:0] mult_wire334 = coe_dat_wire334[9:0] * in_dat_hld334[9:0] ;
    wire [19:0] mult_wire335 = coe_dat_wire335[9:0] * in_dat_hld335[9:0] ;
    wire [19:0] mult_wire336 = coe_dat_wire336[9:0] * in_dat_hld336[9:0] ;
    wire [19:0] mult_wire337 = coe_dat_wire337[9:0] * in_dat_hld337[9:0] ;
    wire [19:0] mult_wire338 = coe_dat_wire338[9:0] * in_dat_hld338[9:0] ;
    wire [19:0] mult_wire339 = coe_dat_wire339[9:0] * in_dat_hld339[9:0] ;
    wire [19:0] mult_wire340 = coe_dat_wire340[9:0] * in_dat_hld340[9:0] ;
    wire [19:0] mult_wire341 = coe_dat_wire341[9:0] * in_dat_hld341[9:0] ;
    wire [19:0] mult_wire342 = coe_dat_wire342[9:0] * in_dat_hld342[9:0] ;
    wire [19:0] mult_wire343 = coe_dat_wire343[9:0] * in_dat_hld343[9:0] ;
    wire [19:0] mult_wire344 = coe_dat_wire344[9:0] * in_dat_hld344[9:0] ;
    wire [19:0] mult_wire345 = coe_dat_wire345[9:0] * in_dat_hld345[9:0] ;
    wire [19:0] mult_wire346 = coe_dat_wire346[9:0] * in_dat_hld346[9:0] ;
    wire [19:0] mult_wire347 = coe_dat_wire347[9:0] * in_dat_hld347[9:0] ;
    wire [19:0] mult_wire348 = coe_dat_wire348[9:0] * in_dat_hld348[9:0] ;
    wire [19:0] mult_wire349 = coe_dat_wire349[9:0] * in_dat_hld349[9:0] ;
    wire [19:0] mult_wire350 = coe_dat_wire350[9:0] * in_dat_hld350[9:0] ;
    wire [19:0] mult_wire351 = coe_dat_wire351[9:0] * in_dat_hld351[9:0] ;
    wire [19:0] mult_wire352 = coe_dat_wire352[9:0] * in_dat_hld352[9:0] ;
    wire [19:0] mult_wire353 = coe_dat_wire353[9:0] * in_dat_hld353[9:0] ;
    wire [19:0] mult_wire354 = coe_dat_wire354[9:0] * in_dat_hld354[9:0] ;
    wire [19:0] mult_wire355 = coe_dat_wire355[9:0] * in_dat_hld355[9:0] ;
    wire [19:0] mult_wire356 = coe_dat_wire356[9:0] * in_dat_hld356[9:0] ;
    wire [19:0] mult_wire357 = coe_dat_wire357[9:0] * in_dat_hld357[9:0] ;
    wire [19:0] mult_wire358 = coe_dat_wire358[9:0] * in_dat_hld358[9:0] ;
    wire [19:0] mult_wire359 = coe_dat_wire359[9:0] * in_dat_hld359[9:0] ;
    wire [19:0] mult_wire360 = coe_dat_wire360[9:0] * in_dat_hld360[9:0] ;
    wire [19:0] mult_wire361 = coe_dat_wire361[9:0] * in_dat_hld361[9:0] ;
    wire [19:0] mult_wire362 = coe_dat_wire362[9:0] * in_dat_hld362[9:0] ;
    wire [19:0] mult_wire363 = coe_dat_wire363[9:0] * in_dat_hld363[9:0] ;
    wire [19:0] mult_wire364 = coe_dat_wire364[9:0] * in_dat_hld364[9:0] ;
    wire [19:0] mult_wire365 = coe_dat_wire365[9:0] * in_dat_hld365[9:0] ;
    wire [19:0] mult_wire366 = coe_dat_wire366[9:0] * in_dat_hld366[9:0] ;
    wire [19:0] mult_wire367 = coe_dat_wire367[9:0] * in_dat_hld367[9:0] ;
    wire [19:0] mult_wire368 = coe_dat_wire368[9:0] * in_dat_hld368[9:0] ;
    wire [19:0] mult_wire369 = coe_dat_wire369[9:0] * in_dat_hld369[9:0] ;
    wire [19:0] mult_wire370 = coe_dat_wire370[9:0] * in_dat_hld370[9:0] ;
    wire [19:0] mult_wire371 = coe_dat_wire371[9:0] * in_dat_hld371[9:0] ;
    wire [19:0] mult_wire372 = coe_dat_wire372[9:0] * in_dat_hld372[9:0] ;
    wire [19:0] mult_wire373 = coe_dat_wire373[9:0] * in_dat_hld373[9:0] ;
    wire [19:0] mult_wire374 = coe_dat_wire374[9:0] * in_dat_hld374[9:0] ;
    wire [19:0] mult_wire375 = coe_dat_wire375[9:0] * in_dat_hld375[9:0] ;
    wire [19:0] mult_wire376 = coe_dat_wire376[9:0] * in_dat_hld376[9:0] ;
    wire [19:0] mult_wire377 = coe_dat_wire377[9:0] * in_dat_hld377[9:0] ;
    wire [19:0] mult_wire378 = coe_dat_wire378[9:0] * in_dat_hld378[9:0] ;
    wire [19:0] mult_wire379 = coe_dat_wire379[9:0] * in_dat_hld379[9:0] ;
    wire [19:0] mult_wire380 = coe_dat_wire380[9:0] * in_dat_hld380[9:0] ;
    wire [19:0] mult_wire381 = coe_dat_wire381[9:0] * in_dat_hld381[9:0] ;
    wire [19:0] mult_wire382 = coe_dat_wire382[9:0] * in_dat_hld382[9:0] ;
    wire [19:0] mult_wire383 = coe_dat_wire383[9:0] * in_dat_hld383[9:0] ;
    wire [19:0] mult_wire384 = coe_dat_wire384[9:0] * in_dat_hld384[9:0] ;
    wire [19:0] mult_wire385 = coe_dat_wire385[9:0] * in_dat_hld385[9:0] ;
    wire [19:0] mult_wire386 = coe_dat_wire386[9:0] * in_dat_hld386[9:0] ;
    wire [19:0] mult_wire387 = coe_dat_wire387[9:0] * in_dat_hld387[9:0] ;
    wire [19:0] mult_wire388 = coe_dat_wire388[9:0] * in_dat_hld388[9:0] ;
    wire [19:0] mult_wire389 = coe_dat_wire389[9:0] * in_dat_hld389[9:0] ;
    wire [19:0] mult_wire390 = coe_dat_wire390[9:0] * in_dat_hld390[9:0] ;
    wire [19:0] mult_wire391 = coe_dat_wire391[9:0] * in_dat_hld391[9:0] ;
    wire [19:0] mult_wire392 = coe_dat_wire392[9:0] * in_dat_hld392[9:0] ;
    wire [19:0] mult_wire393 = coe_dat_wire393[9:0] * in_dat_hld393[9:0] ;
    wire [19:0] mult_wire394 = coe_dat_wire394[9:0] * in_dat_hld394[9:0] ;
    wire [19:0] mult_wire395 = coe_dat_wire395[9:0] * in_dat_hld395[9:0] ;
    wire [19:0] mult_wire396 = coe_dat_wire396[9:0] * in_dat_hld396[9:0] ;
    wire [19:0] mult_wire397 = coe_dat_wire397[9:0] * in_dat_hld397[9:0] ;
    wire [19:0] mult_wire398 = coe_dat_wire398[9:0] * in_dat_hld398[9:0] ;
    wire [19:0] mult_wire399 = coe_dat_wire399[9:0] * in_dat_hld399[9:0] ;
    wire [19:0] mult_wire400 = coe_dat_wire400[9:0] * in_dat_hld400[9:0] ;
    wire [19:0] mult_wire401 = coe_dat_wire401[9:0] * in_dat_hld401[9:0] ;
    wire [19:0] mult_wire402 = coe_dat_wire402[9:0] * in_dat_hld402[9:0] ;
    wire [19:0] mult_wire403 = coe_dat_wire403[9:0] * in_dat_hld403[9:0] ;
    wire [19:0] mult_wire404 = coe_dat_wire404[9:0] * in_dat_hld404[9:0] ;
    wire [19:0] mult_wire405 = coe_dat_wire405[9:0] * in_dat_hld405[9:0] ;
    wire [19:0] mult_wire406 = coe_dat_wire406[9:0] * in_dat_hld406[9:0] ;
    wire [19:0] mult_wire407 = coe_dat_wire407[9:0] * in_dat_hld407[9:0] ;
    wire [19:0] mult_wire408 = coe_dat_wire408[9:0] * in_dat_hld408[9:0] ;
    wire [19:0] mult_wire409 = coe_dat_wire409[9:0] * in_dat_hld409[9:0] ;
    wire [19:0] mult_wire410 = coe_dat_wire410[9:0] * in_dat_hld410[9:0] ;
    wire [19:0] mult_wire411 = coe_dat_wire411[9:0] * in_dat_hld411[9:0] ;
    wire [19:0] mult_wire412 = coe_dat_wire412[9:0] * in_dat_hld412[9:0] ;
    wire [19:0] mult_wire413 = coe_dat_wire413[9:0] * in_dat_hld413[9:0] ;
    wire [19:0] mult_wire414 = coe_dat_wire414[9:0] * in_dat_hld414[9:0] ;
    wire [19:0] mult_wire415 = coe_dat_wire415[9:0] * in_dat_hld415[9:0] ;
    wire [19:0] mult_wire416 = coe_dat_wire416[9:0] * in_dat_hld416[9:0] ;
    wire [19:0] mult_wire417 = coe_dat_wire417[9:0] * in_dat_hld417[9:0] ;
    wire [19:0] mult_wire418 = coe_dat_wire418[9:0] * in_dat_hld418[9:0] ;
    wire [19:0] mult_wire419 = coe_dat_wire419[9:0] * in_dat_hld419[9:0] ;
    wire [19:0] mult_wire420 = coe_dat_wire420[9:0] * in_dat_hld420[9:0] ;
    wire [19:0] mult_wire421 = coe_dat_wire421[9:0] * in_dat_hld421[9:0] ;
    wire [19:0] mult_wire422 = coe_dat_wire422[9:0] * in_dat_hld422[9:0] ;
    wire [19:0] mult_wire423 = coe_dat_wire423[9:0] * in_dat_hld423[9:0] ;
    wire [19:0] mult_wire424 = coe_dat_wire424[9:0] * in_dat_hld424[9:0] ;
    wire [19:0] mult_wire425 = coe_dat_wire425[9:0] * in_dat_hld425[9:0] ;
    wire [19:0] mult_wire426 = coe_dat_wire426[9:0] * in_dat_hld426[9:0] ;
    wire [19:0] mult_wire427 = coe_dat_wire427[9:0] * in_dat_hld427[9:0] ;
    wire [19:0] mult_wire428 = coe_dat_wire428[9:0] * in_dat_hld428[9:0] ;
    wire [19:0] mult_wire429 = coe_dat_wire429[9:0] * in_dat_hld429[9:0] ;
    wire [19:0] mult_wire430 = coe_dat_wire430[9:0] * in_dat_hld430[9:0] ;
    wire [19:0] mult_wire431 = coe_dat_wire431[9:0] * in_dat_hld431[9:0] ;
    wire [19:0] mult_wire432 = coe_dat_wire432[9:0] * in_dat_hld432[9:0] ;
    wire [19:0] mult_wire433 = coe_dat_wire433[9:0] * in_dat_hld433[9:0] ;
    wire [19:0] mult_wire434 = coe_dat_wire434[9:0] * in_dat_hld434[9:0] ;
    wire [19:0] mult_wire435 = coe_dat_wire435[9:0] * in_dat_hld435[9:0] ;
    wire [19:0] mult_wire436 = coe_dat_wire436[9:0] * in_dat_hld436[9:0] ;
    wire [19:0] mult_wire437 = coe_dat_wire437[9:0] * in_dat_hld437[9:0] ;
    wire [19:0] mult_wire438 = coe_dat_wire438[9:0] * in_dat_hld438[9:0] ;
    wire [19:0] mult_wire439 = coe_dat_wire439[9:0] * in_dat_hld439[9:0] ;
    wire [19:0] mult_wire440 = coe_dat_wire440[9:0] * in_dat_hld440[9:0] ;
    wire [19:0] mult_wire441 = coe_dat_wire441[9:0] * in_dat_hld441[9:0] ;
    wire [19:0] mult_wire442 = coe_dat_wire442[9:0] * in_dat_hld442[9:0] ;
    wire [19:0] mult_wire443 = coe_dat_wire443[9:0] * in_dat_hld443[9:0] ;
    wire [19:0] mult_wire444 = coe_dat_wire444[9:0] * in_dat_hld444[9:0] ;
    wire [19:0] mult_wire445 = coe_dat_wire445[9:0] * in_dat_hld445[9:0] ;
    wire [19:0] mult_wire446 = coe_dat_wire446[9:0] * in_dat_hld446[9:0] ;
    wire [19:0] mult_wire447 = coe_dat_wire447[9:0] * in_dat_hld447[9:0] ;
    wire [19:0] mult_wire448 = coe_dat_wire448[9:0] * in_dat_hld448[9:0] ;
    wire [19:0] mult_wire449 = coe_dat_wire449[9:0] * in_dat_hld449[9:0] ;
    wire [19:0] mult_wire450 = coe_dat_wire450[9:0] * in_dat_hld450[9:0] ;
    wire [19:0] mult_wire451 = coe_dat_wire451[9:0] * in_dat_hld451[9:0] ;
    wire [19:0] mult_wire452 = coe_dat_wire452[9:0] * in_dat_hld452[9:0] ;
    wire [19:0] mult_wire453 = coe_dat_wire453[9:0] * in_dat_hld453[9:0] ;
    wire [19:0] mult_wire454 = coe_dat_wire454[9:0] * in_dat_hld454[9:0] ;
    wire [19:0] mult_wire455 = coe_dat_wire455[9:0] * in_dat_hld455[9:0] ;
    wire [19:0] mult_wire456 = coe_dat_wire456[9:0] * in_dat_hld456[9:0] ;
    wire [19:0] mult_wire457 = coe_dat_wire457[9:0] * in_dat_hld457[9:0] ;
    wire [19:0] mult_wire458 = coe_dat_wire458[9:0] * in_dat_hld458[9:0] ;
    wire [19:0] mult_wire459 = coe_dat_wire459[9:0] * in_dat_hld459[9:0] ;
    wire [19:0] mult_wire460 = coe_dat_wire460[9:0] * in_dat_hld460[9:0] ;
    wire [19:0] mult_wire461 = coe_dat_wire461[9:0] * in_dat_hld461[9:0] ;
    wire [19:0] mult_wire462 = coe_dat_wire462[9:0] * in_dat_hld462[9:0] ;
    wire [19:0] mult_wire463 = coe_dat_wire463[9:0] * in_dat_hld463[9:0] ;
    wire [19:0] mult_wire464 = coe_dat_wire464[9:0] * in_dat_hld464[9:0] ;
    wire [19:0] mult_wire465 = coe_dat_wire465[9:0] * in_dat_hld465[9:0] ;
    wire [19:0] mult_wire466 = coe_dat_wire466[9:0] * in_dat_hld466[9:0] ;
    wire [19:0] mult_wire467 = coe_dat_wire467[9:0] * in_dat_hld467[9:0] ;
    wire [19:0] mult_wire468 = coe_dat_wire468[9:0] * in_dat_hld468[9:0] ;
    wire [19:0] mult_wire469 = coe_dat_wire469[9:0] * in_dat_hld469[9:0] ;
    wire [19:0] mult_wire470 = coe_dat_wire470[9:0] * in_dat_hld470[9:0] ;
    wire [19:0] mult_wire471 = coe_dat_wire471[9:0] * in_dat_hld471[9:0] ;
    wire [19:0] mult_wire472 = coe_dat_wire472[9:0] * in_dat_hld472[9:0] ;
    wire [19:0] mult_wire473 = coe_dat_wire473[9:0] * in_dat_hld473[9:0] ;
    wire [19:0] mult_wire474 = coe_dat_wire474[9:0] * in_dat_hld474[9:0] ;
    wire [19:0] mult_wire475 = coe_dat_wire475[9:0] * in_dat_hld475[9:0] ;
    wire [19:0] mult_wire476 = coe_dat_wire476[9:0] * in_dat_hld476[9:0] ;
    wire [19:0] mult_wire477 = coe_dat_wire477[9:0] * in_dat_hld477[9:0] ;
    wire [19:0] mult_wire478 = coe_dat_wire478[9:0] * in_dat_hld478[9:0] ;
    wire [19:0] mult_wire479 = coe_dat_wire479[9:0] * in_dat_hld479[9:0] ;
    wire [19:0] mult_wire480 = coe_dat_wire480[9:0] * in_dat_hld480[9:0] ;
    wire [19:0] mult_wire481 = coe_dat_wire481[9:0] * in_dat_hld481[9:0] ;
    wire [19:0] mult_wire482 = coe_dat_wire482[9:0] * in_dat_hld482[9:0] ;
    wire [19:0] mult_wire483 = coe_dat_wire483[9:0] * in_dat_hld483[9:0] ;
    wire [19:0] mult_wire484 = coe_dat_wire484[9:0] * in_dat_hld484[9:0] ;
    wire [19:0] mult_wire485 = coe_dat_wire485[9:0] * in_dat_hld485[9:0] ;
    wire [19:0] mult_wire486 = coe_dat_wire486[9:0] * in_dat_hld486[9:0] ;
    wire [19:0] mult_wire487 = coe_dat_wire487[9:0] * in_dat_hld487[9:0] ;
    wire [19:0] mult_wire488 = coe_dat_wire488[9:0] * in_dat_hld488[9:0] ;
    wire [19:0] mult_wire489 = coe_dat_wire489[9:0] * in_dat_hld489[9:0] ;
    wire [19:0] mult_wire490 = coe_dat_wire490[9:0] * in_dat_hld490[9:0] ;
    wire [19:0] mult_wire491 = coe_dat_wire491[9:0] * in_dat_hld491[9:0] ;
    wire [19:0] mult_wire492 = coe_dat_wire492[9:0] * in_dat_hld492[9:0] ;
    wire [19:0] mult_wire493 = coe_dat_wire493[9:0] * in_dat_hld493[9:0] ;
    wire [19:0] mult_wire494 = coe_dat_wire494[9:0] * in_dat_hld494[9:0] ;
    wire [19:0] mult_wire495 = coe_dat_wire495[9:0] * in_dat_hld495[9:0] ;
    wire [19:0] mult_wire496 = coe_dat_wire496[9:0] * in_dat_hld496[9:0] ;
    wire [19:0] mult_wire497 = coe_dat_wire497[9:0] * in_dat_hld497[9:0] ;
    wire [19:0] mult_wire498 = coe_dat_wire498[9:0] * in_dat_hld498[9:0] ;
    wire [19:0] mult_wire499 = coe_dat_wire499[9:0] * in_dat_hld499[9:0] ;
    wire [19:0] mult_wire500 = coe_dat_wire500[9:0] * in_dat_hld500[9:0] ;
    wire [19:0] mult_wire501 = coe_dat_wire501[9:0] * in_dat_hld501[9:0] ;
    wire [19:0] mult_wire502 = coe_dat_wire502[9:0] * in_dat_hld502[9:0] ;
    wire [19:0] mult_wire503 = coe_dat_wire503[9:0] * in_dat_hld503[9:0] ;
    wire [19:0] mult_wire504 = coe_dat_wire504[9:0] * in_dat_hld504[9:0] ;
    wire [19:0] mult_wire505 = coe_dat_wire505[9:0] * in_dat_hld505[9:0] ;
    wire [19:0] mult_wire506 = coe_dat_wire506[9:0] * in_dat_hld506[9:0] ;
    wire [19:0] mult_wire507 = coe_dat_wire507[9:0] * in_dat_hld507[9:0] ;
    wire [19:0] mult_wire508 = coe_dat_wire508[9:0] * in_dat_hld508[9:0] ;
    wire [19:0] mult_wire509 = coe_dat_wire509[9:0] * in_dat_hld509[9:0] ;
    wire [19:0] mult_wire510 = coe_dat_wire510[9:0] * in_dat_hld510[9:0] ;
    wire [19:0] mult_wire511 = coe_dat_wire511[9:0] * in_dat_hld511[9:0] ;
    wire [19:0] mult_wire512 = coe_dat_wire512[9:0] * in_dat_hld512[9:0] ;
//
    reg [19:0] mult_reg01,  mult_reg02,  mult_reg03,  mult_reg04,
               mult_reg05,  mult_reg06,  mult_reg07,  mult_reg08,
               mult_reg09,  mult_reg10,  mult_reg11,  mult_reg12,
               mult_reg13,  mult_reg14,  mult_reg15,  mult_reg16,
               mult_reg17,  mult_reg18,  mult_reg19,  mult_reg20,
               mult_reg21,  mult_reg22,  mult_reg23,  mult_reg24,
               mult_reg25,  mult_reg26,  mult_reg27,  mult_reg28,
               mult_reg29,  mult_reg30,  mult_reg31,  mult_reg32,
               mult_reg33,  mult_reg34,  mult_reg35,  mult_reg36,
               mult_reg37,  mult_reg38,  mult_reg39,  mult_reg40,
               mult_reg41,  mult_reg42,  mult_reg43,  mult_reg44,
               mult_reg45,  mult_reg46,  mult_reg47,  mult_reg48,
               mult_reg49,  mult_reg50,  mult_reg51,  mult_reg52,
               mult_reg53,  mult_reg54,  mult_reg55,  mult_reg56,
               mult_reg57,  mult_reg58,  mult_reg59,  mult_reg60,
               mult_reg61,  mult_reg62,  mult_reg63,  mult_reg64,
               mult_reg65,  mult_reg66,  mult_reg67,  mult_reg68,
               mult_reg69,  mult_reg70,  mult_reg71,  mult_reg72,
               mult_reg73,  mult_reg74,  mult_reg75,  mult_reg76,
               mult_reg77,  mult_reg78,  mult_reg79,  mult_reg80,
               mult_reg81,  mult_reg82,  mult_reg83,  mult_reg84,
               mult_reg85,  mult_reg86,  mult_reg87,  mult_reg88,
               mult_reg89,  mult_reg90,  mult_reg91,  mult_reg92,
               mult_reg93,  mult_reg94,  mult_reg95,  mult_reg96,
               mult_reg97,  mult_reg98,  mult_reg99,  mult_reg100,
               mult_reg101, mult_reg102, mult_reg103, mult_reg104,
               mult_reg105, mult_reg106, mult_reg107, mult_reg108,
               mult_reg109, mult_reg110, mult_reg111, mult_reg112,
               mult_reg113, mult_reg114, mult_reg115, mult_reg116,
               mult_reg117, mult_reg118, mult_reg119, mult_reg120,
               mult_reg121, mult_reg122, mult_reg123, mult_reg124,
               mult_reg125, mult_reg126, mult_reg127, mult_reg128,
               mult_reg129, mult_reg130, mult_reg131, mult_reg132,
               mult_reg133, mult_reg134, mult_reg135, mult_reg136,
               mult_reg137, mult_reg138, mult_reg139, mult_reg140,
               mult_reg141, mult_reg142, mult_reg143, mult_reg144,
               mult_reg145, mult_reg146, mult_reg147, mult_reg148,
               mult_reg149, mult_reg150, mult_reg151, mult_reg152,
               mult_reg153, mult_reg154, mult_reg155, mult_reg156,
               mult_reg157, mult_reg158, mult_reg159, mult_reg160,
               mult_reg161, mult_reg162, mult_reg163, mult_reg164,
               mult_reg165, mult_reg166, mult_reg167, mult_reg168,
               mult_reg169, mult_reg170, mult_reg171, mult_reg172,
               mult_reg173, mult_reg174, mult_reg175, mult_reg176,
               mult_reg177, mult_reg178, mult_reg179, mult_reg180,
               mult_reg181, mult_reg182, mult_reg183, mult_reg184,
               mult_reg185, mult_reg186, mult_reg187, mult_reg188,
               mult_reg189, mult_reg190, mult_reg191, mult_reg192,
               mult_reg193, mult_reg194, mult_reg195, mult_reg196,
               mult_reg197, mult_reg198, mult_reg199, mult_reg200,
               mult_reg201, mult_reg202, mult_reg203, mult_reg204,
               mult_reg205, mult_reg206, mult_reg207, mult_reg208,
               mult_reg209, mult_reg210, mult_reg211, mult_reg212,
               mult_reg213, mult_reg214, mult_reg215, mult_reg216,
               mult_reg217, mult_reg218, mult_reg219, mult_reg220,
               mult_reg221, mult_reg222, mult_reg223, mult_reg224,
               mult_reg225, mult_reg226, mult_reg227, mult_reg228,
               mult_reg229, mult_reg230, mult_reg231, mult_reg232,
               mult_reg233, mult_reg234, mult_reg235, mult_reg236,
               mult_reg237, mult_reg238, mult_reg239, mult_reg240,
               mult_reg241, mult_reg242, mult_reg243, mult_reg244,
               mult_reg245, mult_reg246, mult_reg247, mult_reg248,
               mult_reg249, mult_reg250, mult_reg251, mult_reg252,
               mult_reg253, mult_reg254, mult_reg255, mult_reg256,
               mult_reg257, mult_reg258, mult_reg259, mult_reg260,
               mult_reg261, mult_reg262, mult_reg263, mult_reg264,
               mult_reg265, mult_reg266, mult_reg267, mult_reg268,
               mult_reg269, mult_reg270, mult_reg271, mult_reg272,
               mult_reg273, mult_reg274, mult_reg275, mult_reg276,
               mult_reg277, mult_reg278, mult_reg279, mult_reg280,
               mult_reg281, mult_reg282, mult_reg283, mult_reg284,
               mult_reg285, mult_reg286, mult_reg287, mult_reg288,
               mult_reg289, mult_reg290, mult_reg291, mult_reg292,
               mult_reg293, mult_reg294, mult_reg295, mult_reg296,
               mult_reg297, mult_reg298, mult_reg299, mult_reg300,
               mult_reg301, mult_reg302, mult_reg303, mult_reg304,
               mult_reg305, mult_reg306, mult_reg307, mult_reg308,
               mult_reg309, mult_reg310, mult_reg311, mult_reg312,
               mult_reg313, mult_reg314, mult_reg315, mult_reg316,
               mult_reg317, mult_reg318, mult_reg319, mult_reg320,
               mult_reg321, mult_reg322, mult_reg323, mult_reg324,
               mult_reg325, mult_reg326, mult_reg327, mult_reg328,
               mult_reg329, mult_reg330, mult_reg331, mult_reg332,
               mult_reg333, mult_reg334, mult_reg335, mult_reg336,
               mult_reg337, mult_reg338, mult_reg339, mult_reg340,
               mult_reg341, mult_reg342, mult_reg343, mult_reg344,
               mult_reg345, mult_reg346, mult_reg347, mult_reg348,
               mult_reg349, mult_reg350, mult_reg351, mult_reg352,
               mult_reg353, mult_reg354, mult_reg355, mult_reg356,
               mult_reg357, mult_reg358, mult_reg359, mult_reg360,
               mult_reg361, mult_reg362, mult_reg363, mult_reg364,
               mult_reg365, mult_reg366, mult_reg367, mult_reg368,
               mult_reg369, mult_reg370, mult_reg371, mult_reg372,
               mult_reg373, mult_reg374, mult_reg375, mult_reg376,
               mult_reg377, mult_reg378, mult_reg379, mult_reg380,
               mult_reg381, mult_reg382, mult_reg383, mult_reg384,
               mult_reg385, mult_reg386, mult_reg387, mult_reg388,
               mult_reg389, mult_reg390, mult_reg391, mult_reg392,
               mult_reg393, mult_reg394, mult_reg395, mult_reg396,
               mult_reg397, mult_reg398, mult_reg399, mult_reg400,
               mult_reg401, mult_reg402, mult_reg403, mult_reg404,
               mult_reg405, mult_reg406, mult_reg407, mult_reg408,
               mult_reg409, mult_reg410, mult_reg411, mult_reg412,
               mult_reg413, mult_reg414, mult_reg415, mult_reg416,
               mult_reg417, mult_reg418, mult_reg419, mult_reg420,
               mult_reg421, mult_reg422, mult_reg423, mult_reg424,
               mult_reg425, mult_reg426, mult_reg427, mult_reg428,
               mult_reg429, mult_reg430, mult_reg431, mult_reg432,
               mult_reg433, mult_reg434, mult_reg435, mult_reg436,
               mult_reg437, mult_reg438, mult_reg439, mult_reg440,
               mult_reg441, mult_reg442, mult_reg443, mult_reg444,
               mult_reg445, mult_reg446, mult_reg447, mult_reg448,
               mult_reg449, mult_reg450, mult_reg451, mult_reg452,
               mult_reg453, mult_reg454, mult_reg455, mult_reg456,
               mult_reg457, mult_reg458, mult_reg459, mult_reg460,
               mult_reg461, mult_reg462, mult_reg463, mult_reg464,
               mult_reg465, mult_reg466, mult_reg467, mult_reg468,
               mult_reg469, mult_reg470, mult_reg471, mult_reg472,
               mult_reg473, mult_reg474, mult_reg475, mult_reg476,
               mult_reg477, mult_reg478, mult_reg479, mult_reg480,
               mult_reg481, mult_reg482, mult_reg483, mult_reg484,
               mult_reg485, mult_reg486, mult_reg487, mult_reg488,
               mult_reg489, mult_reg490, mult_reg491, mult_reg492,
               mult_reg493, mult_reg494, mult_reg495, mult_reg496,
               mult_reg497, mult_reg498, mult_reg499, mult_reg500,
               mult_reg501, mult_reg502, mult_reg503, mult_reg504,
               mult_reg505, mult_reg506, mult_reg507, mult_reg508,
               mult_reg509, mult_reg510, mult_reg511, mult_reg512;


    always @ (posedge clk) begin
		if(rst) begin
            mult_reg01[19:0]  <= #DLY 20'd0 ;
            mult_reg02[19:0]  <= #DLY 20'd0 ;
            mult_reg03[19:0]  <= #DLY 20'd0 ;
            mult_reg04[19:0]  <= #DLY 20'd0 ;
            mult_reg05[19:0]  <= #DLY 20'd0 ;
            mult_reg06[19:0]  <= #DLY 20'd0 ;
            mult_reg07[19:0]  <= #DLY 20'd0 ;
            mult_reg08[19:0]  <= #DLY 20'd0 ;
            mult_reg09[19:0]  <= #DLY 20'd0 ;
            mult_reg10[19:0]  <= #DLY 20'd0 ;
            mult_reg11[19:0]  <= #DLY 20'd0 ;
            mult_reg12[19:0]  <= #DLY 20'd0 ;
            mult_reg13[19:0]  <= #DLY 20'd0 ;
            mult_reg14[19:0]  <= #DLY 20'd0 ;
            mult_reg15[19:0]  <= #DLY 20'd0 ;
            mult_reg16[19:0]  <= #DLY 20'd0 ;
            mult_reg17[19:0]  <= #DLY 20'd0 ;
            mult_reg18[19:0]  <= #DLY 20'd0 ;
            mult_reg19[19:0]  <= #DLY 20'd0 ;
            mult_reg20[19:0]  <= #DLY 20'd0 ;
            mult_reg21[19:0]  <= #DLY 20'd0 ;
            mult_reg22[19:0]  <= #DLY 20'd0 ;
            mult_reg23[19:0]  <= #DLY 20'd0 ;
            mult_reg24[19:0]  <= #DLY 20'd0 ;
            mult_reg25[19:0]  <= #DLY 20'd0 ;
            mult_reg26[19:0]  <= #DLY 20'd0 ;
            mult_reg27[19:0]  <= #DLY 20'd0 ;
            mult_reg28[19:0]  <= #DLY 20'd0 ;
            mult_reg29[19:0]  <= #DLY 20'd0 ;
            mult_reg30[19:0]  <= #DLY 20'd0 ;
            mult_reg31[19:0]  <= #DLY 20'd0 ;
            mult_reg32[19:0]  <= #DLY 20'd0 ;
            mult_reg33[19:0]  <= #DLY 20'd0 ;
            mult_reg34[19:0]  <= #DLY 20'd0 ;
            mult_reg35[19:0]  <= #DLY 20'd0 ;
            mult_reg36[19:0]  <= #DLY 20'd0 ;
            mult_reg37[19:0]  <= #DLY 20'd0 ;
            mult_reg38[19:0]  <= #DLY 20'd0 ;
            mult_reg39[19:0]  <= #DLY 20'd0 ;
            mult_reg40[19:0]  <= #DLY 20'd0 ;
            mult_reg41[19:0]  <= #DLY 20'd0 ;
            mult_reg42[19:0]  <= #DLY 20'd0 ;
            mult_reg43[19:0]  <= #DLY 20'd0 ;
            mult_reg44[19:0]  <= #DLY 20'd0 ;
            mult_reg45[19:0]  <= #DLY 20'd0 ;
            mult_reg46[19:0]  <= #DLY 20'd0 ;
            mult_reg47[19:0]  <= #DLY 20'd0 ;
            mult_reg48[19:0]  <= #DLY 20'd0 ;
            mult_reg49[19:0]  <= #DLY 20'd0 ;
            mult_reg50[19:0]  <= #DLY 20'd0 ;
            mult_reg51[19:0]  <= #DLY 20'd0 ;
            mult_reg52[19:0]  <= #DLY 20'd0 ;
            mult_reg53[19:0]  <= #DLY 20'd0 ;
            mult_reg54[19:0]  <= #DLY 20'd0 ;
            mult_reg55[19:0]  <= #DLY 20'd0 ;
            mult_reg56[19:0]  <= #DLY 20'd0 ;
            mult_reg57[19:0]  <= #DLY 20'd0 ;
            mult_reg58[19:0]  <= #DLY 20'd0 ;
            mult_reg59[19:0]  <= #DLY 20'd0 ;
            mult_reg60[19:0]  <= #DLY 20'd0 ;
            mult_reg61[19:0]  <= #DLY 20'd0 ;
            mult_reg62[19:0]  <= #DLY 20'd0 ;
            mult_reg63[19:0]  <= #DLY 20'd0 ;
            mult_reg64[19:0]  <= #DLY 20'd0 ;
            mult_reg65[19:0]  <= #DLY 20'd0 ;
            mult_reg66[19:0]  <= #DLY 20'd0 ;
            mult_reg67[19:0]  <= #DLY 20'd0 ;
            mult_reg68[19:0]  <= #DLY 20'd0 ;
            mult_reg69[19:0]  <= #DLY 20'd0 ;
            mult_reg70[19:0]  <= #DLY 20'd0 ;
            mult_reg71[19:0]  <= #DLY 20'd0 ;
            mult_reg72[19:0]  <= #DLY 20'd0 ;
            mult_reg73[19:0]  <= #DLY 20'd0 ;
            mult_reg74[19:0]  <= #DLY 20'd0 ;
            mult_reg75[19:0]  <= #DLY 20'd0 ;
            mult_reg76[19:0]  <= #DLY 20'd0 ;
            mult_reg77[19:0]  <= #DLY 20'd0 ;
            mult_reg78[19:0]  <= #DLY 20'd0 ;
            mult_reg79[19:0]  <= #DLY 20'd0 ;
            mult_reg80[19:0]  <= #DLY 20'd0 ;
            mult_reg81[19:0]  <= #DLY 20'd0 ;
            mult_reg82[19:0]  <= #DLY 20'd0 ;
            mult_reg83[19:0]  <= #DLY 20'd0 ;
            mult_reg84[19:0]  <= #DLY 20'd0 ;
            mult_reg85[19:0]  <= #DLY 20'd0 ;
            mult_reg86[19:0]  <= #DLY 20'd0 ;
            mult_reg87[19:0]  <= #DLY 20'd0 ;
            mult_reg88[19:0]  <= #DLY 20'd0 ;
            mult_reg89[19:0]  <= #DLY 20'd0 ;
            mult_reg90[19:0]  <= #DLY 20'd0 ;
            mult_reg91[19:0]  <= #DLY 20'd0 ;
            mult_reg92[19:0]  <= #DLY 20'd0 ;
            mult_reg93[19:0]  <= #DLY 20'd0 ;
            mult_reg94[19:0]  <= #DLY 20'd0 ;
            mult_reg95[19:0]  <= #DLY 20'd0 ;
            mult_reg96[19:0]  <= #DLY 20'd0 ;
            mult_reg97[19:0]  <= #DLY 20'd0 ;
            mult_reg98[19:0]  <= #DLY 20'd0 ;
            mult_reg99[19:0]  <= #DLY 20'd0 ;
            mult_reg100[19:0] <= #DLY 20'd0 ;
            mult_reg101[19:0] <= #DLY 20'd0 ;
            mult_reg102[19:0] <= #DLY 20'd0 ;
            mult_reg103[19:0] <= #DLY 20'd0 ;
            mult_reg104[19:0] <= #DLY 20'd0 ;
            mult_reg105[19:0] <= #DLY 20'd0 ;
            mult_reg106[19:0] <= #DLY 20'd0 ;
            mult_reg107[19:0] <= #DLY 20'd0 ;
            mult_reg108[19:0] <= #DLY 20'd0 ;
            mult_reg109[19:0] <= #DLY 20'd0 ;
            mult_reg110[19:0] <= #DLY 20'd0 ;
            mult_reg111[19:0] <= #DLY 20'd0 ;
            mult_reg112[19:0] <= #DLY 20'd0 ;
            mult_reg113[19:0] <= #DLY 20'd0 ;
            mult_reg114[19:0] <= #DLY 20'd0 ;
            mult_reg115[19:0] <= #DLY 20'd0 ;
            mult_reg116[19:0] <= #DLY 20'd0 ;
            mult_reg117[19:0] <= #DLY 20'd0 ;
            mult_reg118[19:0] <= #DLY 20'd0 ;
            mult_reg119[19:0] <= #DLY 20'd0 ;
            mult_reg120[19:0] <= #DLY 20'd0 ;
            mult_reg121[19:0] <= #DLY 20'd0 ;
            mult_reg122[19:0] <= #DLY 20'd0 ;
            mult_reg123[19:0] <= #DLY 20'd0 ;
            mult_reg124[19:0] <= #DLY 20'd0 ;
            mult_reg125[19:0] <= #DLY 20'd0 ;
            mult_reg126[19:0] <= #DLY 20'd0 ;
            mult_reg127[19:0] <= #DLY 20'd0 ;
            mult_reg128[19:0] <= #DLY 20'd0 ;
            mult_reg129[19:0] <= #DLY 20'd0 ;
            mult_reg130[19:0] <= #DLY 20'd0 ;
            mult_reg131[19:0] <= #DLY 20'd0 ;
            mult_reg132[19:0] <= #DLY 20'd0 ;
            mult_reg133[19:0] <= #DLY 20'd0 ;
            mult_reg134[19:0] <= #DLY 20'd0 ;
            mult_reg135[19:0] <= #DLY 20'd0 ;
            mult_reg136[19:0] <= #DLY 20'd0 ;
            mult_reg137[19:0] <= #DLY 20'd0 ;
            mult_reg138[19:0] <= #DLY 20'd0 ;
            mult_reg139[19:0] <= #DLY 20'd0 ;
            mult_reg140[19:0] <= #DLY 20'd0 ;
            mult_reg141[19:0] <= #DLY 20'd0 ;
            mult_reg142[19:0] <= #DLY 20'd0 ;
            mult_reg143[19:0] <= #DLY 20'd0 ;
            mult_reg144[19:0] <= #DLY 20'd0 ;
            mult_reg145[19:0] <= #DLY 20'd0 ;
            mult_reg146[19:0] <= #DLY 20'd0 ;
            mult_reg147[19:0] <= #DLY 20'd0 ;
            mult_reg148[19:0] <= #DLY 20'd0 ;
            mult_reg149[19:0] <= #DLY 20'd0 ;
            mult_reg150[19:0] <= #DLY 20'd0 ;
            mult_reg151[19:0] <= #DLY 20'd0 ;
            mult_reg152[19:0] <= #DLY 20'd0 ;
            mult_reg153[19:0] <= #DLY 20'd0 ;
            mult_reg154[19:0] <= #DLY 20'd0 ;
            mult_reg155[19:0] <= #DLY 20'd0 ;
            mult_reg156[19:0] <= #DLY 20'd0 ;
            mult_reg157[19:0] <= #DLY 20'd0 ;
            mult_reg158[19:0] <= #DLY 20'd0 ;
            mult_reg159[19:0] <= #DLY 20'd0 ;
            mult_reg160[19:0] <= #DLY 20'd0 ;
            mult_reg161[19:0] <= #DLY 20'd0 ;
            mult_reg162[19:0] <= #DLY 20'd0 ;
            mult_reg163[19:0] <= #DLY 20'd0 ;
            mult_reg164[19:0] <= #DLY 20'd0 ;
            mult_reg165[19:0] <= #DLY 20'd0 ;
            mult_reg166[19:0] <= #DLY 20'd0 ;
            mult_reg167[19:0] <= #DLY 20'd0 ;
            mult_reg168[19:0] <= #DLY 20'd0 ;
            mult_reg169[19:0] <= #DLY 20'd0 ;
            mult_reg170[19:0] <= #DLY 20'd0 ;
            mult_reg171[19:0] <= #DLY 20'd0 ;
            mult_reg172[19:0] <= #DLY 20'd0 ;
            mult_reg173[19:0] <= #DLY 20'd0 ;
            mult_reg174[19:0] <= #DLY 20'd0 ;
            mult_reg175[19:0] <= #DLY 20'd0 ;
            mult_reg176[19:0] <= #DLY 20'd0 ;
            mult_reg177[19:0] <= #DLY 20'd0 ;
            mult_reg178[19:0] <= #DLY 20'd0 ;
            mult_reg179[19:0] <= #DLY 20'd0 ;
            mult_reg180[19:0] <= #DLY 20'd0 ;
            mult_reg181[19:0] <= #DLY 20'd0 ;
            mult_reg182[19:0] <= #DLY 20'd0 ;
            mult_reg183[19:0] <= #DLY 20'd0 ;
            mult_reg184[19:0] <= #DLY 20'd0 ;
            mult_reg185[19:0] <= #DLY 20'd0 ;
            mult_reg186[19:0] <= #DLY 20'd0 ;
            mult_reg187[19:0] <= #DLY 20'd0 ;
            mult_reg188[19:0] <= #DLY 20'd0 ;
            mult_reg189[19:0] <= #DLY 20'd0 ;
            mult_reg190[19:0] <= #DLY 20'd0 ;
            mult_reg191[19:0] <= #DLY 20'd0 ;
            mult_reg192[19:0] <= #DLY 20'd0 ;
            mult_reg193[19:0] <= #DLY 20'd0 ;
            mult_reg194[19:0] <= #DLY 20'd0 ;
            mult_reg195[19:0] <= #DLY 20'd0 ;
            mult_reg196[19:0] <= #DLY 20'd0 ;
            mult_reg197[19:0] <= #DLY 20'd0 ;
            mult_reg198[19:0] <= #DLY 20'd0 ;
            mult_reg199[19:0] <= #DLY 20'd0 ;
            mult_reg200[19:0] <= #DLY 20'd0 ;
            mult_reg201[19:0] <= #DLY 20'd0 ;
            mult_reg202[19:0] <= #DLY 20'd0 ;
            mult_reg203[19:0] <= #DLY 20'd0 ;
            mult_reg204[19:0] <= #DLY 20'd0 ;
            mult_reg205[19:0] <= #DLY 20'd0 ;
            mult_reg206[19:0] <= #DLY 20'd0 ;
            mult_reg207[19:0] <= #DLY 20'd0 ;
            mult_reg208[19:0] <= #DLY 20'd0 ;
            mult_reg209[19:0] <= #DLY 20'd0 ;
            mult_reg210[19:0] <= #DLY 20'd0 ;
            mult_reg211[19:0] <= #DLY 20'd0 ;
            mult_reg212[19:0] <= #DLY 20'd0 ;
            mult_reg213[19:0] <= #DLY 20'd0 ;
            mult_reg214[19:0] <= #DLY 20'd0 ;
            mult_reg215[19:0] <= #DLY 20'd0 ;
            mult_reg216[19:0] <= #DLY 20'd0 ;
            mult_reg217[19:0] <= #DLY 20'd0 ;
            mult_reg218[19:0] <= #DLY 20'd0 ;
            mult_reg219[19:0] <= #DLY 20'd0 ;
            mult_reg220[19:0] <= #DLY 20'd0 ;
            mult_reg221[19:0] <= #DLY 20'd0 ;
            mult_reg222[19:0] <= #DLY 20'd0 ;
            mult_reg223[19:0] <= #DLY 20'd0 ;
            mult_reg224[19:0] <= #DLY 20'd0 ;
            mult_reg225[19:0] <= #DLY 20'd0 ;
            mult_reg226[19:0] <= #DLY 20'd0 ;
            mult_reg227[19:0] <= #DLY 20'd0 ;
            mult_reg228[19:0] <= #DLY 20'd0 ;
            mult_reg229[19:0] <= #DLY 20'd0 ;
            mult_reg230[19:0] <= #DLY 20'd0 ;
            mult_reg231[19:0] <= #DLY 20'd0 ;
            mult_reg232[19:0] <= #DLY 20'd0 ;
            mult_reg233[19:0] <= #DLY 20'd0 ;
            mult_reg234[19:0] <= #DLY 20'd0 ;
            mult_reg235[19:0] <= #DLY 20'd0 ;
            mult_reg236[19:0] <= #DLY 20'd0 ;
            mult_reg237[19:0] <= #DLY 20'd0 ;
            mult_reg238[19:0] <= #DLY 20'd0 ;
            mult_reg239[19:0] <= #DLY 20'd0 ;
            mult_reg240[19:0] <= #DLY 20'd0 ;
            mult_reg241[19:0] <= #DLY 20'd0 ;
            mult_reg242[19:0] <= #DLY 20'd0 ;
            mult_reg243[19:0] <= #DLY 20'd0 ;
            mult_reg244[19:0] <= #DLY 20'd0 ;
            mult_reg245[19:0] <= #DLY 20'd0 ;
            mult_reg246[19:0] <= #DLY 20'd0 ;
            mult_reg247[19:0] <= #DLY 20'd0 ;
            mult_reg248[19:0] <= #DLY 20'd0 ;
            mult_reg249[19:0] <= #DLY 20'd0 ;
            mult_reg250[19:0] <= #DLY 20'd0 ;
            mult_reg251[19:0] <= #DLY 20'd0 ;
            mult_reg252[19:0] <= #DLY 20'd0 ;
            mult_reg253[19:0] <= #DLY 20'd0 ;
            mult_reg254[19:0] <= #DLY 20'd0 ;
            mult_reg255[19:0] <= #DLY 20'd0 ;
            mult_reg256[19:0] <= #DLY 20'd0 ;
            mult_reg257[19:0] <= #DLY 20'd0 ;
            mult_reg258[19:0] <= #DLY 20'd0 ;
            mult_reg259[19:0] <= #DLY 20'd0 ;
            mult_reg260[19:0] <= #DLY 20'd0 ;
            mult_reg261[19:0] <= #DLY 20'd0 ;
            mult_reg262[19:0] <= #DLY 20'd0 ;
            mult_reg263[19:0] <= #DLY 20'd0 ;
            mult_reg264[19:0] <= #DLY 20'd0 ;
            mult_reg265[19:0] <= #DLY 20'd0 ;
            mult_reg266[19:0] <= #DLY 20'd0 ;
            mult_reg267[19:0] <= #DLY 20'd0 ;
            mult_reg268[19:0] <= #DLY 20'd0 ;
            mult_reg269[19:0] <= #DLY 20'd0 ;
            mult_reg270[19:0] <= #DLY 20'd0 ;
            mult_reg271[19:0] <= #DLY 20'd0 ;
            mult_reg272[19:0] <= #DLY 20'd0 ;
            mult_reg273[19:0] <= #DLY 20'd0 ;
            mult_reg274[19:0] <= #DLY 20'd0 ;
            mult_reg275[19:0] <= #DLY 20'd0 ;
            mult_reg276[19:0] <= #DLY 20'd0 ;
            mult_reg277[19:0] <= #DLY 20'd0 ;
            mult_reg278[19:0] <= #DLY 20'd0 ;
            mult_reg279[19:0] <= #DLY 20'd0 ;
            mult_reg280[19:0] <= #DLY 20'd0 ;
            mult_reg281[19:0] <= #DLY 20'd0 ;
            mult_reg282[19:0] <= #DLY 20'd0 ;
            mult_reg283[19:0] <= #DLY 20'd0 ;
            mult_reg284[19:0] <= #DLY 20'd0 ;
            mult_reg285[19:0] <= #DLY 20'd0 ;
            mult_reg286[19:0] <= #DLY 20'd0 ;
            mult_reg287[19:0] <= #DLY 20'd0 ;
            mult_reg288[19:0] <= #DLY 20'd0 ;
            mult_reg289[19:0] <= #DLY 20'd0 ;
            mult_reg290[19:0] <= #DLY 20'd0 ;
            mult_reg291[19:0] <= #DLY 20'd0 ;
            mult_reg292[19:0] <= #DLY 20'd0 ;
            mult_reg293[19:0] <= #DLY 20'd0 ;
            mult_reg294[19:0] <= #DLY 20'd0 ;
            mult_reg295[19:0] <= #DLY 20'd0 ;
            mult_reg296[19:0] <= #DLY 20'd0 ;
            mult_reg297[19:0] <= #DLY 20'd0 ;
            mult_reg298[19:0] <= #DLY 20'd0 ;
            mult_reg299[19:0] <= #DLY 20'd0 ;
            mult_reg300[19:0] <= #DLY 20'd0 ;
            mult_reg301[19:0] <= #DLY 20'd0 ;
            mult_reg302[19:0] <= #DLY 20'd0 ;
            mult_reg303[19:0] <= #DLY 20'd0 ;
            mult_reg304[19:0] <= #DLY 20'd0 ;
            mult_reg305[19:0] <= #DLY 20'd0 ;
            mult_reg306[19:0] <= #DLY 20'd0 ;
            mult_reg307[19:0] <= #DLY 20'd0 ;
            mult_reg308[19:0] <= #DLY 20'd0 ;
            mult_reg309[19:0] <= #DLY 20'd0 ;
            mult_reg310[19:0] <= #DLY 20'd0 ;
            mult_reg311[19:0] <= #DLY 20'd0 ;
            mult_reg312[19:0] <= #DLY 20'd0 ;
            mult_reg313[19:0] <= #DLY 20'd0 ;
            mult_reg314[19:0] <= #DLY 20'd0 ;
            mult_reg315[19:0] <= #DLY 20'd0 ;
            mult_reg316[19:0] <= #DLY 20'd0 ;
            mult_reg317[19:0] <= #DLY 20'd0 ;
            mult_reg318[19:0] <= #DLY 20'd0 ;
            mult_reg319[19:0] <= #DLY 20'd0 ;
            mult_reg320[19:0] <= #DLY 20'd0 ;
            mult_reg321[19:0] <= #DLY 20'd0 ;
            mult_reg322[19:0] <= #DLY 20'd0 ;
            mult_reg323[19:0] <= #DLY 20'd0 ;
            mult_reg324[19:0] <= #DLY 20'd0 ;
            mult_reg325[19:0] <= #DLY 20'd0 ;
            mult_reg326[19:0] <= #DLY 20'd0 ;
            mult_reg327[19:0] <= #DLY 20'd0 ;
            mult_reg328[19:0] <= #DLY 20'd0 ;
            mult_reg329[19:0] <= #DLY 20'd0 ;
            mult_reg330[19:0] <= #DLY 20'd0 ;
            mult_reg331[19:0] <= #DLY 20'd0 ;
            mult_reg332[19:0] <= #DLY 20'd0 ;
            mult_reg333[19:0] <= #DLY 20'd0 ;
            mult_reg334[19:0] <= #DLY 20'd0 ;
            mult_reg335[19:0] <= #DLY 20'd0 ;
            mult_reg336[19:0] <= #DLY 20'd0 ;
            mult_reg337[19:0] <= #DLY 20'd0 ;
            mult_reg338[19:0] <= #DLY 20'd0 ;
            mult_reg339[19:0] <= #DLY 20'd0 ;
            mult_reg340[19:0] <= #DLY 20'd0 ;
            mult_reg341[19:0] <= #DLY 20'd0 ;
            mult_reg342[19:0] <= #DLY 20'd0 ;
            mult_reg343[19:0] <= #DLY 20'd0 ;
            mult_reg344[19:0] <= #DLY 20'd0 ;
            mult_reg345[19:0] <= #DLY 20'd0 ;
            mult_reg346[19:0] <= #DLY 20'd0 ;
            mult_reg347[19:0] <= #DLY 20'd0 ;
            mult_reg348[19:0] <= #DLY 20'd0 ;
            mult_reg349[19:0] <= #DLY 20'd0 ;
            mult_reg350[19:0] <= #DLY 20'd0 ;
            mult_reg351[19:0] <= #DLY 20'd0 ;
            mult_reg352[19:0] <= #DLY 20'd0 ;
            mult_reg353[19:0] <= #DLY 20'd0 ;
            mult_reg354[19:0] <= #DLY 20'd0 ;
            mult_reg355[19:0] <= #DLY 20'd0 ;
            mult_reg356[19:0] <= #DLY 20'd0 ;
            mult_reg357[19:0] <= #DLY 20'd0 ;
            mult_reg358[19:0] <= #DLY 20'd0 ;
            mult_reg359[19:0] <= #DLY 20'd0 ;
            mult_reg360[19:0] <= #DLY 20'd0 ;
            mult_reg361[19:0] <= #DLY 20'd0 ;
            mult_reg362[19:0] <= #DLY 20'd0 ;
            mult_reg363[19:0] <= #DLY 20'd0 ;
            mult_reg364[19:0] <= #DLY 20'd0 ;
            mult_reg365[19:0] <= #DLY 20'd0 ;
            mult_reg366[19:0] <= #DLY 20'd0 ;
            mult_reg367[19:0] <= #DLY 20'd0 ;
            mult_reg368[19:0] <= #DLY 20'd0 ;
            mult_reg369[19:0] <= #DLY 20'd0 ;
            mult_reg370[19:0] <= #DLY 20'd0 ;
            mult_reg371[19:0] <= #DLY 20'd0 ;
            mult_reg372[19:0] <= #DLY 20'd0 ;
            mult_reg373[19:0] <= #DLY 20'd0 ;
            mult_reg374[19:0] <= #DLY 20'd0 ;
            mult_reg375[19:0] <= #DLY 20'd0 ;
            mult_reg376[19:0] <= #DLY 20'd0 ;
            mult_reg377[19:0] <= #DLY 20'd0 ;
            mult_reg378[19:0] <= #DLY 20'd0 ;
            mult_reg379[19:0] <= #DLY 20'd0 ;
            mult_reg380[19:0] <= #DLY 20'd0 ;
            mult_reg381[19:0] <= #DLY 20'd0 ;
            mult_reg382[19:0] <= #DLY 20'd0 ;
            mult_reg383[19:0] <= #DLY 20'd0 ;
            mult_reg384[19:0] <= #DLY 20'd0 ;
            mult_reg385[19:0] <= #DLY 20'd0 ;
            mult_reg386[19:0] <= #DLY 20'd0 ;
            mult_reg387[19:0] <= #DLY 20'd0 ;
            mult_reg388[19:0] <= #DLY 20'd0 ;
            mult_reg389[19:0] <= #DLY 20'd0 ;
            mult_reg390[19:0] <= #DLY 20'd0 ;
            mult_reg391[19:0] <= #DLY 20'd0 ;
            mult_reg392[19:0] <= #DLY 20'd0 ;
            mult_reg393[19:0] <= #DLY 20'd0 ;
            mult_reg394[19:0] <= #DLY 20'd0 ;
            mult_reg395[19:0] <= #DLY 20'd0 ;
            mult_reg396[19:0] <= #DLY 20'd0 ;
            mult_reg397[19:0] <= #DLY 20'd0 ;
            mult_reg398[19:0] <= #DLY 20'd0 ;
            mult_reg399[19:0] <= #DLY 20'd0 ;
            mult_reg400[19:0] <= #DLY 20'd0 ;
            mult_reg401[19:0] <= #DLY 20'd0 ;
            mult_reg402[19:0] <= #DLY 20'd0 ;
            mult_reg403[19:0] <= #DLY 20'd0 ;
            mult_reg404[19:0] <= #DLY 20'd0 ;
            mult_reg405[19:0] <= #DLY 20'd0 ;
            mult_reg406[19:0] <= #DLY 20'd0 ;
            mult_reg407[19:0] <= #DLY 20'd0 ;
            mult_reg408[19:0] <= #DLY 20'd0 ;
            mult_reg409[19:0] <= #DLY 20'd0 ;
            mult_reg410[19:0] <= #DLY 20'd0 ;
            mult_reg411[19:0] <= #DLY 20'd0 ;
            mult_reg412[19:0] <= #DLY 20'd0 ;
            mult_reg413[19:0] <= #DLY 20'd0 ;
            mult_reg414[19:0] <= #DLY 20'd0 ;
            mult_reg415[19:0] <= #DLY 20'd0 ;
            mult_reg416[19:0] <= #DLY 20'd0 ;
            mult_reg417[19:0] <= #DLY 20'd0 ;
            mult_reg418[19:0] <= #DLY 20'd0 ;
            mult_reg419[19:0] <= #DLY 20'd0 ;
            mult_reg420[19:0] <= #DLY 20'd0 ;
            mult_reg421[19:0] <= #DLY 20'd0 ;
            mult_reg422[19:0] <= #DLY 20'd0 ;
            mult_reg423[19:0] <= #DLY 20'd0 ;
            mult_reg424[19:0] <= #DLY 20'd0 ;
            mult_reg425[19:0] <= #DLY 20'd0 ;
            mult_reg426[19:0] <= #DLY 20'd0 ;
            mult_reg427[19:0] <= #DLY 20'd0 ;
            mult_reg428[19:0] <= #DLY 20'd0 ;
            mult_reg429[19:0] <= #DLY 20'd0 ;
            mult_reg430[19:0] <= #DLY 20'd0 ;
            mult_reg431[19:0] <= #DLY 20'd0 ;
            mult_reg432[19:0] <= #DLY 20'd0 ;
            mult_reg433[19:0] <= #DLY 20'd0 ;
            mult_reg434[19:0] <= #DLY 20'd0 ;
            mult_reg435[19:0] <= #DLY 20'd0 ;
            mult_reg436[19:0] <= #DLY 20'd0 ;
            mult_reg437[19:0] <= #DLY 20'd0 ;
            mult_reg438[19:0] <= #DLY 20'd0 ;
            mult_reg439[19:0] <= #DLY 20'd0 ;
            mult_reg440[19:0] <= #DLY 20'd0 ;
            mult_reg441[19:0] <= #DLY 20'd0 ;
            mult_reg442[19:0] <= #DLY 20'd0 ;
            mult_reg443[19:0] <= #DLY 20'd0 ;
            mult_reg444[19:0] <= #DLY 20'd0 ;
            mult_reg445[19:0] <= #DLY 20'd0 ;
            mult_reg446[19:0] <= #DLY 20'd0 ;
            mult_reg447[19:0] <= #DLY 20'd0 ;
            mult_reg448[19:0] <= #DLY 20'd0 ;
            mult_reg449[19:0] <= #DLY 20'd0 ;
            mult_reg450[19:0] <= #DLY 20'd0 ;
            mult_reg451[19:0] <= #DLY 20'd0 ;
            mult_reg452[19:0] <= #DLY 20'd0 ;
            mult_reg453[19:0] <= #DLY 20'd0 ;
            mult_reg454[19:0] <= #DLY 20'd0 ;
            mult_reg455[19:0] <= #DLY 20'd0 ;
            mult_reg456[19:0] <= #DLY 20'd0 ;
            mult_reg457[19:0] <= #DLY 20'd0 ;
            mult_reg458[19:0] <= #DLY 20'd0 ;
            mult_reg459[19:0] <= #DLY 20'd0 ;
            mult_reg460[19:0] <= #DLY 20'd0 ;
            mult_reg461[19:0] <= #DLY 20'd0 ;
            mult_reg462[19:0] <= #DLY 20'd0 ;
            mult_reg463[19:0] <= #DLY 20'd0 ;
            mult_reg464[19:0] <= #DLY 20'd0 ;
            mult_reg465[19:0] <= #DLY 20'd0 ;
            mult_reg466[19:0] <= #DLY 20'd0 ;
            mult_reg467[19:0] <= #DLY 20'd0 ;
            mult_reg468[19:0] <= #DLY 20'd0 ;
            mult_reg469[19:0] <= #DLY 20'd0 ;
            mult_reg470[19:0] <= #DLY 20'd0 ;
            mult_reg471[19:0] <= #DLY 20'd0 ;
            mult_reg472[19:0] <= #DLY 20'd0 ;
            mult_reg473[19:0] <= #DLY 20'd0 ;
            mult_reg474[19:0] <= #DLY 20'd0 ;
            mult_reg475[19:0] <= #DLY 20'd0 ;
            mult_reg476[19:0] <= #DLY 20'd0 ;
            mult_reg477[19:0] <= #DLY 20'd0 ;
            mult_reg478[19:0] <= #DLY 20'd0 ;
            mult_reg479[19:0] <= #DLY 20'd0 ;
            mult_reg480[19:0] <= #DLY 20'd0 ;
            mult_reg481[19:0] <= #DLY 20'd0 ;
            mult_reg482[19:0] <= #DLY 20'd0 ;
            mult_reg483[19:0] <= #DLY 20'd0 ;
            mult_reg484[19:0] <= #DLY 20'd0 ;
            mult_reg485[19:0] <= #DLY 20'd0 ;
            mult_reg486[19:0] <= #DLY 20'd0 ;
            mult_reg487[19:0] <= #DLY 20'd0 ;
            mult_reg488[19:0] <= #DLY 20'd0 ;
            mult_reg489[19:0] <= #DLY 20'd0 ;
            mult_reg490[19:0] <= #DLY 20'd0 ;
            mult_reg491[19:0] <= #DLY 20'd0 ;
            mult_reg492[19:0] <= #DLY 20'd0 ;
            mult_reg493[19:0] <= #DLY 20'd0 ;
            mult_reg494[19:0] <= #DLY 20'd0 ;
            mult_reg495[19:0] <= #DLY 20'd0 ;
            mult_reg496[19:0] <= #DLY 20'd0 ;
            mult_reg497[19:0] <= #DLY 20'd0 ;
            mult_reg498[19:0] <= #DLY 20'd0 ;
            mult_reg499[19:0] <= #DLY 20'd0 ;
            mult_reg500[19:0] <= #DLY 20'd0 ;
            mult_reg501[19:0] <= #DLY 20'd0 ;
            mult_reg502[19:0] <= #DLY 20'd0 ;
            mult_reg503[19:0] <= #DLY 20'd0 ;
            mult_reg504[19:0] <= #DLY 20'd0 ;
            mult_reg505[19:0] <= #DLY 20'd0 ;
            mult_reg506[19:0] <= #DLY 20'd0 ;
            mult_reg507[19:0] <= #DLY 20'd0 ;
            mult_reg508[19:0] <= #DLY 20'd0 ;
            mult_reg509[19:0] <= #DLY 20'd0 ;
            mult_reg510[19:0] <= #DLY 20'd0 ;
            mult_reg511[19:0] <= #DLY 20'd0 ;
            mult_reg512[19:0] <= #DLY 20'd0 ;
		end else begin
            mult_reg01[19:0]  <= #DLY mult_wire01[19:0]  ;
            mult_reg02[19:0]  <= #DLY mult_wire02[19:0]  ;
            mult_reg03[19:0]  <= #DLY mult_wire03[19:0]  ;
            mult_reg04[19:0]  <= #DLY mult_wire04[19:0]  ;
            mult_reg05[19:0]  <= #DLY mult_wire05[19:0]  ;
            mult_reg06[19:0]  <= #DLY mult_wire06[19:0]  ;
            mult_reg07[19:0]  <= #DLY mult_wire07[19:0]  ;
            mult_reg08[19:0]  <= #DLY mult_wire08[19:0]  ;
            mult_reg09[19:0]  <= #DLY mult_wire09[19:0]  ;
            mult_reg10[19:0]  <= #DLY mult_wire10[19:0]  ;
            mult_reg11[19:0]  <= #DLY mult_wire11[19:0]  ;
            mult_reg12[19:0]  <= #DLY mult_wire12[19:0]  ;
            mult_reg13[19:0]  <= #DLY mult_wire13[19:0]  ;
            mult_reg14[19:0]  <= #DLY mult_wire14[19:0]  ;
            mult_reg15[19:0]  <= #DLY mult_wire15[19:0]  ;
            mult_reg16[19:0]  <= #DLY mult_wire16[19:0]  ;
            mult_reg17[19:0]  <= #DLY mult_wire17[19:0]  ;
            mult_reg18[19:0]  <= #DLY mult_wire18[19:0]  ;
            mult_reg19[19:0]  <= #DLY mult_wire19[19:0]  ;
            mult_reg20[19:0]  <= #DLY mult_wire20[19:0]  ;
            mult_reg21[19:0]  <= #DLY mult_wire21[19:0]  ;
            mult_reg22[19:0]  <= #DLY mult_wire22[19:0]  ;
            mult_reg23[19:0]  <= #DLY mult_wire23[19:0]  ;
            mult_reg24[19:0]  <= #DLY mult_wire24[19:0]  ;
            mult_reg25[19:0]  <= #DLY mult_wire25[19:0]  ;
            mult_reg26[19:0]  <= #DLY mult_wire26[19:0]  ;
            mult_reg27[19:0]  <= #DLY mult_wire27[19:0]  ;
            mult_reg28[19:0]  <= #DLY mult_wire28[19:0]  ;
            mult_reg29[19:0]  <= #DLY mult_wire29[19:0]  ;
            mult_reg30[19:0]  <= #DLY mult_wire30[19:0]  ;
            mult_reg31[19:0]  <= #DLY mult_wire31[19:0]  ;
            mult_reg32[19:0]  <= #DLY mult_wire32[19:0]  ;
            mult_reg33[19:0]  <= #DLY mult_wire33[19:0]  ;
            mult_reg34[19:0]  <= #DLY mult_wire34[19:0]  ;
            mult_reg35[19:0]  <= #DLY mult_wire35[19:0]  ;
            mult_reg36[19:0]  <= #DLY mult_wire36[19:0]  ;
            mult_reg37[19:0]  <= #DLY mult_wire37[19:0]  ;
            mult_reg38[19:0]  <= #DLY mult_wire38[19:0]  ;
            mult_reg39[19:0]  <= #DLY mult_wire39[19:0]  ;
            mult_reg40[19:0]  <= #DLY mult_wire40[19:0]  ;
            mult_reg41[19:0]  <= #DLY mult_wire41[19:0]  ;
            mult_reg42[19:0]  <= #DLY mult_wire42[19:0]  ;
            mult_reg43[19:0]  <= #DLY mult_wire43[19:0]  ;
            mult_reg44[19:0]  <= #DLY mult_wire44[19:0]  ;
            mult_reg45[19:0]  <= #DLY mult_wire45[19:0]  ;
            mult_reg46[19:0]  <= #DLY mult_wire46[19:0]  ;
            mult_reg47[19:0]  <= #DLY mult_wire47[19:0]  ;
            mult_reg48[19:0]  <= #DLY mult_wire48[19:0]  ;
            mult_reg49[19:0]  <= #DLY mult_wire49[19:0]  ;
            mult_reg50[19:0]  <= #DLY mult_wire50[19:0]  ;
            mult_reg51[19:0]  <= #DLY mult_wire51[19:0]  ;
            mult_reg52[19:0]  <= #DLY mult_wire52[19:0]  ;
            mult_reg53[19:0]  <= #DLY mult_wire53[19:0]  ;
            mult_reg54[19:0]  <= #DLY mult_wire54[19:0]  ;
            mult_reg55[19:0]  <= #DLY mult_wire55[19:0]  ;
            mult_reg56[19:0]  <= #DLY mult_wire56[19:0]  ;
            mult_reg57[19:0]  <= #DLY mult_wire57[19:0]  ;
            mult_reg58[19:0]  <= #DLY mult_wire58[19:0]  ;
            mult_reg59[19:0]  <= #DLY mult_wire59[19:0]  ;
            mult_reg60[19:0]  <= #DLY mult_wire60[19:0]  ;
            mult_reg61[19:0]  <= #DLY mult_wire61[19:0]  ;
            mult_reg62[19:0]  <= #DLY mult_wire62[19:0]  ;
            mult_reg63[19:0]  <= #DLY mult_wire63[19:0]  ;
            mult_reg64[19:0]  <= #DLY mult_wire64[19:0]  ;
            mult_reg65[19:0]  <= #DLY mult_wire65[19:0]  ;
            mult_reg66[19:0]  <= #DLY mult_wire66[19:0]  ;
            mult_reg67[19:0]  <= #DLY mult_wire67[19:0]  ;
            mult_reg68[19:0]  <= #DLY mult_wire68[19:0]  ;
            mult_reg69[19:0]  <= #DLY mult_wire69[19:0]  ;
            mult_reg70[19:0]  <= #DLY mult_wire70[19:0]  ;
            mult_reg71[19:0]  <= #DLY mult_wire71[19:0]  ;
            mult_reg72[19:0]  <= #DLY mult_wire72[19:0]  ;
            mult_reg73[19:0]  <= #DLY mult_wire73[19:0]  ;
            mult_reg74[19:0]  <= #DLY mult_wire74[19:0]  ;
            mult_reg75[19:0]  <= #DLY mult_wire75[19:0]  ;
            mult_reg76[19:0]  <= #DLY mult_wire76[19:0]  ;
            mult_reg77[19:0]  <= #DLY mult_wire77[19:0]  ;
            mult_reg78[19:0]  <= #DLY mult_wire78[19:0]  ;
            mult_reg79[19:0]  <= #DLY mult_wire79[19:0]  ;
            mult_reg80[19:0]  <= #DLY mult_wire80[19:0]  ;
            mult_reg81[19:0]  <= #DLY mult_wire81[19:0]  ;
            mult_reg82[19:0]  <= #DLY mult_wire82[19:0]  ;
            mult_reg83[19:0]  <= #DLY mult_wire83[19:0]  ;
            mult_reg84[19:0]  <= #DLY mult_wire84[19:0]  ;
            mult_reg85[19:0]  <= #DLY mult_wire85[19:0]  ;
            mult_reg86[19:0]  <= #DLY mult_wire86[19:0]  ;
            mult_reg87[19:0]  <= #DLY mult_wire87[19:0]  ;
            mult_reg88[19:0]  <= #DLY mult_wire88[19:0]  ;
            mult_reg89[19:0]  <= #DLY mult_wire89[19:0]  ;
            mult_reg90[19:0]  <= #DLY mult_wire90[19:0]  ;
            mult_reg91[19:0]  <= #DLY mult_wire91[19:0]  ;
            mult_reg92[19:0]  <= #DLY mult_wire92[19:0]  ;
            mult_reg93[19:0]  <= #DLY mult_wire93[19:0]  ;
            mult_reg94[19:0]  <= #DLY mult_wire94[19:0]  ;
            mult_reg95[19:0]  <= #DLY mult_wire95[19:0]  ;
            mult_reg96[19:0]  <= #DLY mult_wire96[19:0]  ;
            mult_reg97[19:0]  <= #DLY mult_wire97[19:0]  ;
            mult_reg98[19:0]  <= #DLY mult_wire98[19:0]  ;
            mult_reg99[19:0]  <= #DLY mult_wire99[19:0]  ;
            mult_reg100[19:0] <= #DLY mult_wire100[19:0] ;
            mult_reg101[19:0] <= #DLY mult_wire101[19:0] ;
            mult_reg102[19:0] <= #DLY mult_wire102[19:0] ;
            mult_reg103[19:0] <= #DLY mult_wire103[19:0] ;
            mult_reg104[19:0] <= #DLY mult_wire104[19:0] ;
            mult_reg105[19:0] <= #DLY mult_wire105[19:0] ;
            mult_reg106[19:0] <= #DLY mult_wire106[19:0] ;
            mult_reg107[19:0] <= #DLY mult_wire107[19:0] ;
            mult_reg108[19:0] <= #DLY mult_wire108[19:0] ;
            mult_reg109[19:0] <= #DLY mult_wire109[19:0] ;
            mult_reg110[19:0] <= #DLY mult_wire110[19:0] ;
            mult_reg111[19:0] <= #DLY mult_wire111[19:0] ;
            mult_reg112[19:0] <= #DLY mult_wire112[19:0] ;
            mult_reg113[19:0] <= #DLY mult_wire113[19:0] ;
            mult_reg114[19:0] <= #DLY mult_wire114[19:0] ;
            mult_reg115[19:0] <= #DLY mult_wire115[19:0] ;
            mult_reg116[19:0] <= #DLY mult_wire116[19:0] ;
            mult_reg117[19:0] <= #DLY mult_wire117[19:0] ;
            mult_reg118[19:0] <= #DLY mult_wire118[19:0] ;
            mult_reg119[19:0] <= #DLY mult_wire119[19:0] ;
            mult_reg120[19:0] <= #DLY mult_wire120[19:0] ;
            mult_reg121[19:0] <= #DLY mult_wire121[19:0] ;
            mult_reg122[19:0] <= #DLY mult_wire122[19:0] ;
            mult_reg123[19:0] <= #DLY mult_wire123[19:0] ;
            mult_reg124[19:0] <= #DLY mult_wire124[19:0] ;
            mult_reg125[19:0] <= #DLY mult_wire125[19:0] ;
            mult_reg126[19:0] <= #DLY mult_wire126[19:0] ;
            mult_reg127[19:0] <= #DLY mult_wire127[19:0] ;
            mult_reg128[19:0] <= #DLY mult_wire128[19:0] ;
            mult_reg129[19:0] <= #DLY mult_wire129[19:0] ;
            mult_reg130[19:0] <= #DLY mult_wire130[19:0] ;
            mult_reg131[19:0] <= #DLY mult_wire131[19:0] ;
            mult_reg132[19:0] <= #DLY mult_wire132[19:0] ;
            mult_reg133[19:0] <= #DLY mult_wire133[19:0] ;
            mult_reg134[19:0] <= #DLY mult_wire134[19:0] ;
            mult_reg135[19:0] <= #DLY mult_wire135[19:0] ;
            mult_reg136[19:0] <= #DLY mult_wire136[19:0] ;
            mult_reg137[19:0] <= #DLY mult_wire137[19:0] ;
            mult_reg138[19:0] <= #DLY mult_wire138[19:0] ;
            mult_reg139[19:0] <= #DLY mult_wire139[19:0] ;
            mult_reg140[19:0] <= #DLY mult_wire140[19:0] ;
            mult_reg141[19:0] <= #DLY mult_wire141[19:0] ;
            mult_reg142[19:0] <= #DLY mult_wire142[19:0] ;
            mult_reg143[19:0] <= #DLY mult_wire143[19:0] ;
            mult_reg144[19:0] <= #DLY mult_wire144[19:0] ;
            mult_reg145[19:0] <= #DLY mult_wire145[19:0] ;
            mult_reg146[19:0] <= #DLY mult_wire146[19:0] ;
            mult_reg147[19:0] <= #DLY mult_wire147[19:0] ;
            mult_reg148[19:0] <= #DLY mult_wire148[19:0] ;
            mult_reg149[19:0] <= #DLY mult_wire149[19:0] ;
            mult_reg150[19:0] <= #DLY mult_wire150[19:0] ;
            mult_reg151[19:0] <= #DLY mult_wire151[19:0] ;
            mult_reg152[19:0] <= #DLY mult_wire152[19:0] ;
            mult_reg153[19:0] <= #DLY mult_wire153[19:0] ;
            mult_reg154[19:0] <= #DLY mult_wire154[19:0] ;
            mult_reg155[19:0] <= #DLY mult_wire155[19:0] ;
            mult_reg156[19:0] <= #DLY mult_wire156[19:0] ;
            mult_reg157[19:0] <= #DLY mult_wire157[19:0] ;
            mult_reg158[19:0] <= #DLY mult_wire158[19:0] ;
            mult_reg159[19:0] <= #DLY mult_wire159[19:0] ;
            mult_reg160[19:0] <= #DLY mult_wire160[19:0] ;
            mult_reg161[19:0] <= #DLY mult_wire161[19:0] ;
            mult_reg162[19:0] <= #DLY mult_wire162[19:0] ;
            mult_reg163[19:0] <= #DLY mult_wire163[19:0] ;
            mult_reg164[19:0] <= #DLY mult_wire164[19:0] ;
            mult_reg165[19:0] <= #DLY mult_wire165[19:0] ;
            mult_reg166[19:0] <= #DLY mult_wire166[19:0] ;
            mult_reg167[19:0] <= #DLY mult_wire167[19:0] ;
            mult_reg168[19:0] <= #DLY mult_wire168[19:0] ;
            mult_reg169[19:0] <= #DLY mult_wire169[19:0] ;
            mult_reg170[19:0] <= #DLY mult_wire170[19:0] ;
            mult_reg171[19:0] <= #DLY mult_wire171[19:0] ;
            mult_reg172[19:0] <= #DLY mult_wire172[19:0] ;
            mult_reg173[19:0] <= #DLY mult_wire173[19:0] ;
            mult_reg174[19:0] <= #DLY mult_wire174[19:0] ;
            mult_reg175[19:0] <= #DLY mult_wire175[19:0] ;
            mult_reg176[19:0] <= #DLY mult_wire176[19:0] ;
            mult_reg177[19:0] <= #DLY mult_wire177[19:0] ;
            mult_reg178[19:0] <= #DLY mult_wire178[19:0] ;
            mult_reg179[19:0] <= #DLY mult_wire179[19:0] ;
            mult_reg180[19:0] <= #DLY mult_wire180[19:0] ;
            mult_reg181[19:0] <= #DLY mult_wire181[19:0] ;
            mult_reg182[19:0] <= #DLY mult_wire182[19:0] ;
            mult_reg183[19:0] <= #DLY mult_wire183[19:0] ;
            mult_reg184[19:0] <= #DLY mult_wire184[19:0] ;
            mult_reg185[19:0] <= #DLY mult_wire185[19:0] ;
            mult_reg186[19:0] <= #DLY mult_wire186[19:0] ;
            mult_reg187[19:0] <= #DLY mult_wire187[19:0] ;
            mult_reg188[19:0] <= #DLY mult_wire188[19:0] ;
            mult_reg189[19:0] <= #DLY mult_wire189[19:0] ;
            mult_reg190[19:0] <= #DLY mult_wire190[19:0] ;
            mult_reg191[19:0] <= #DLY mult_wire191[19:0] ;
            mult_reg192[19:0] <= #DLY mult_wire192[19:0] ;
            mult_reg193[19:0] <= #DLY mult_wire193[19:0] ;
            mult_reg194[19:0] <= #DLY mult_wire194[19:0] ;
            mult_reg195[19:0] <= #DLY mult_wire195[19:0] ;
            mult_reg196[19:0] <= #DLY mult_wire196[19:0] ;
            mult_reg197[19:0] <= #DLY mult_wire197[19:0] ;
            mult_reg198[19:0] <= #DLY mult_wire198[19:0] ;
            mult_reg199[19:0] <= #DLY mult_wire199[19:0] ;
            mult_reg200[19:0] <= #DLY mult_wire200[19:0] ;
            mult_reg201[19:0] <= #DLY mult_wire201[19:0] ;
            mult_reg202[19:0] <= #DLY mult_wire202[19:0] ;
            mult_reg203[19:0] <= #DLY mult_wire203[19:0] ;
            mult_reg204[19:0] <= #DLY mult_wire204[19:0] ;
            mult_reg205[19:0] <= #DLY mult_wire205[19:0] ;
            mult_reg206[19:0] <= #DLY mult_wire206[19:0] ;
            mult_reg207[19:0] <= #DLY mult_wire207[19:0] ;
            mult_reg208[19:0] <= #DLY mult_wire208[19:0] ;
            mult_reg209[19:0] <= #DLY mult_wire209[19:0] ;
            mult_reg210[19:0] <= #DLY mult_wire210[19:0] ;
            mult_reg211[19:0] <= #DLY mult_wire211[19:0] ;
            mult_reg212[19:0] <= #DLY mult_wire212[19:0] ;
            mult_reg213[19:0] <= #DLY mult_wire213[19:0] ;
            mult_reg214[19:0] <= #DLY mult_wire214[19:0] ;
            mult_reg215[19:0] <= #DLY mult_wire215[19:0] ;
            mult_reg216[19:0] <= #DLY mult_wire216[19:0] ;
            mult_reg217[19:0] <= #DLY mult_wire217[19:0] ;
            mult_reg218[19:0] <= #DLY mult_wire218[19:0] ;
            mult_reg219[19:0] <= #DLY mult_wire219[19:0] ;
            mult_reg220[19:0] <= #DLY mult_wire220[19:0] ;
            mult_reg221[19:0] <= #DLY mult_wire221[19:0] ;
            mult_reg222[19:0] <= #DLY mult_wire222[19:0] ;
            mult_reg223[19:0] <= #DLY mult_wire223[19:0] ;
            mult_reg224[19:0] <= #DLY mult_wire224[19:0] ;
            mult_reg225[19:0] <= #DLY mult_wire225[19:0] ;
            mult_reg226[19:0] <= #DLY mult_wire226[19:0] ;
            mult_reg227[19:0] <= #DLY mult_wire227[19:0] ;
            mult_reg228[19:0] <= #DLY mult_wire228[19:0] ;
            mult_reg229[19:0] <= #DLY mult_wire229[19:0] ;
            mult_reg230[19:0] <= #DLY mult_wire230[19:0] ;
            mult_reg231[19:0] <= #DLY mult_wire231[19:0] ;
            mult_reg232[19:0] <= #DLY mult_wire232[19:0] ;
            mult_reg233[19:0] <= #DLY mult_wire233[19:0] ;
            mult_reg234[19:0] <= #DLY mult_wire234[19:0] ;
            mult_reg235[19:0] <= #DLY mult_wire235[19:0] ;
            mult_reg236[19:0] <= #DLY mult_wire236[19:0] ;
            mult_reg237[19:0] <= #DLY mult_wire237[19:0] ;
            mult_reg238[19:0] <= #DLY mult_wire238[19:0] ;
            mult_reg239[19:0] <= #DLY mult_wire239[19:0] ;
            mult_reg240[19:0] <= #DLY mult_wire240[19:0] ;
            mult_reg241[19:0] <= #DLY mult_wire241[19:0] ;
            mult_reg242[19:0] <= #DLY mult_wire242[19:0] ;
            mult_reg243[19:0] <= #DLY mult_wire243[19:0] ;
            mult_reg244[19:0] <= #DLY mult_wire244[19:0] ;
            mult_reg245[19:0] <= #DLY mult_wire245[19:0] ;
            mult_reg246[19:0] <= #DLY mult_wire246[19:0] ;
            mult_reg247[19:0] <= #DLY mult_wire247[19:0] ;
            mult_reg248[19:0] <= #DLY mult_wire248[19:0] ;
            mult_reg249[19:0] <= #DLY mult_wire249[19:0] ;
            mult_reg250[19:0] <= #DLY mult_wire250[19:0] ;
            mult_reg251[19:0] <= #DLY mult_wire251[19:0] ;
            mult_reg252[19:0] <= #DLY mult_wire252[19:0] ;
            mult_reg253[19:0] <= #DLY mult_wire253[19:0] ;
            mult_reg254[19:0] <= #DLY mult_wire254[19:0] ;
            mult_reg255[19:0] <= #DLY mult_wire255[19:0] ;
            mult_reg256[19:0] <= #DLY mult_wire256[19:0] ;
            mult_reg257[19:0] <= #DLY mult_wire257[19:0] ;
            mult_reg258[19:0] <= #DLY mult_wire258[19:0] ;
            mult_reg259[19:0] <= #DLY mult_wire259[19:0] ;
            mult_reg260[19:0] <= #DLY mult_wire260[19:0] ;
            mult_reg261[19:0] <= #DLY mult_wire261[19:0] ;
            mult_reg262[19:0] <= #DLY mult_wire262[19:0] ;
            mult_reg263[19:0] <= #DLY mult_wire263[19:0] ;
            mult_reg264[19:0] <= #DLY mult_wire264[19:0] ;
            mult_reg265[19:0] <= #DLY mult_wire265[19:0] ;
            mult_reg266[19:0] <= #DLY mult_wire266[19:0] ;
            mult_reg267[19:0] <= #DLY mult_wire267[19:0] ;
            mult_reg268[19:0] <= #DLY mult_wire268[19:0] ;
            mult_reg269[19:0] <= #DLY mult_wire269[19:0] ;
            mult_reg270[19:0] <= #DLY mult_wire270[19:0] ;
            mult_reg271[19:0] <= #DLY mult_wire271[19:0] ;
            mult_reg272[19:0] <= #DLY mult_wire272[19:0] ;
            mult_reg273[19:0] <= #DLY mult_wire273[19:0] ;
            mult_reg274[19:0] <= #DLY mult_wire274[19:0] ;
            mult_reg275[19:0] <= #DLY mult_wire275[19:0] ;
            mult_reg276[19:0] <= #DLY mult_wire276[19:0] ;
            mult_reg277[19:0] <= #DLY mult_wire277[19:0] ;
            mult_reg278[19:0] <= #DLY mult_wire278[19:0] ;
            mult_reg279[19:0] <= #DLY mult_wire279[19:0] ;
            mult_reg280[19:0] <= #DLY mult_wire280[19:0] ;
            mult_reg281[19:0] <= #DLY mult_wire281[19:0] ;
            mult_reg282[19:0] <= #DLY mult_wire282[19:0] ;
            mult_reg283[19:0] <= #DLY mult_wire283[19:0] ;
            mult_reg284[19:0] <= #DLY mult_wire284[19:0] ;
            mult_reg285[19:0] <= #DLY mult_wire285[19:0] ;
            mult_reg286[19:0] <= #DLY mult_wire286[19:0] ;
            mult_reg287[19:0] <= #DLY mult_wire287[19:0] ;
            mult_reg288[19:0] <= #DLY mult_wire288[19:0] ;
            mult_reg289[19:0] <= #DLY mult_wire289[19:0] ;
            mult_reg290[19:0] <= #DLY mult_wire290[19:0] ;
            mult_reg291[19:0] <= #DLY mult_wire291[19:0] ;
            mult_reg292[19:0] <= #DLY mult_wire292[19:0] ;
            mult_reg293[19:0] <= #DLY mult_wire293[19:0] ;
            mult_reg294[19:0] <= #DLY mult_wire294[19:0] ;
            mult_reg295[19:0] <= #DLY mult_wire295[19:0] ;
            mult_reg296[19:0] <= #DLY mult_wire296[19:0] ;
            mult_reg297[19:0] <= #DLY mult_wire297[19:0] ;
            mult_reg298[19:0] <= #DLY mult_wire298[19:0] ;
            mult_reg299[19:0] <= #DLY mult_wire299[19:0] ;
            mult_reg300[19:0] <= #DLY mult_wire300[19:0] ;
            mult_reg301[19:0] <= #DLY mult_wire301[19:0] ;
            mult_reg302[19:0] <= #DLY mult_wire302[19:0] ;
            mult_reg303[19:0] <= #DLY mult_wire303[19:0] ;
            mult_reg304[19:0] <= #DLY mult_wire304[19:0] ;
            mult_reg305[19:0] <= #DLY mult_wire305[19:0] ;
            mult_reg306[19:0] <= #DLY mult_wire306[19:0] ;
            mult_reg307[19:0] <= #DLY mult_wire307[19:0] ;
            mult_reg308[19:0] <= #DLY mult_wire308[19:0] ;
            mult_reg309[19:0] <= #DLY mult_wire309[19:0] ;
            mult_reg310[19:0] <= #DLY mult_wire310[19:0] ;
            mult_reg311[19:0] <= #DLY mult_wire311[19:0] ;
            mult_reg312[19:0] <= #DLY mult_wire312[19:0] ;
            mult_reg313[19:0] <= #DLY mult_wire313[19:0] ;
            mult_reg314[19:0] <= #DLY mult_wire314[19:0] ;
            mult_reg315[19:0] <= #DLY mult_wire315[19:0] ;
            mult_reg316[19:0] <= #DLY mult_wire316[19:0] ;
            mult_reg317[19:0] <= #DLY mult_wire317[19:0] ;
            mult_reg318[19:0] <= #DLY mult_wire318[19:0] ;
            mult_reg319[19:0] <= #DLY mult_wire319[19:0] ;
            mult_reg320[19:0] <= #DLY mult_wire320[19:0] ;
            mult_reg321[19:0] <= #DLY mult_wire321[19:0] ;
            mult_reg322[19:0] <= #DLY mult_wire322[19:0] ;
            mult_reg323[19:0] <= #DLY mult_wire323[19:0] ;
            mult_reg324[19:0] <= #DLY mult_wire324[19:0] ;
            mult_reg325[19:0] <= #DLY mult_wire325[19:0] ;
            mult_reg326[19:0] <= #DLY mult_wire326[19:0] ;
            mult_reg327[19:0] <= #DLY mult_wire327[19:0] ;
            mult_reg328[19:0] <= #DLY mult_wire328[19:0] ;
            mult_reg329[19:0] <= #DLY mult_wire329[19:0] ;
            mult_reg330[19:0] <= #DLY mult_wire330[19:0] ;
            mult_reg331[19:0] <= #DLY mult_wire331[19:0] ;
            mult_reg332[19:0] <= #DLY mult_wire332[19:0] ;
            mult_reg333[19:0] <= #DLY mult_wire333[19:0] ;
            mult_reg334[19:0] <= #DLY mult_wire334[19:0] ;
            mult_reg335[19:0] <= #DLY mult_wire335[19:0] ;
            mult_reg336[19:0] <= #DLY mult_wire336[19:0] ;
            mult_reg337[19:0] <= #DLY mult_wire337[19:0] ;
            mult_reg338[19:0] <= #DLY mult_wire338[19:0] ;
            mult_reg339[19:0] <= #DLY mult_wire339[19:0] ;
            mult_reg340[19:0] <= #DLY mult_wire340[19:0] ;
            mult_reg341[19:0] <= #DLY mult_wire341[19:0] ;
            mult_reg342[19:0] <= #DLY mult_wire342[19:0] ;
            mult_reg343[19:0] <= #DLY mult_wire343[19:0] ;
            mult_reg344[19:0] <= #DLY mult_wire344[19:0] ;
            mult_reg345[19:0] <= #DLY mult_wire345[19:0] ;
            mult_reg346[19:0] <= #DLY mult_wire346[19:0] ;
            mult_reg347[19:0] <= #DLY mult_wire347[19:0] ;
            mult_reg348[19:0] <= #DLY mult_wire348[19:0] ;
            mult_reg349[19:0] <= #DLY mult_wire349[19:0] ;
            mult_reg350[19:0] <= #DLY mult_wire350[19:0] ;
            mult_reg351[19:0] <= #DLY mult_wire351[19:0] ;
            mult_reg352[19:0] <= #DLY mult_wire352[19:0] ;
            mult_reg353[19:0] <= #DLY mult_wire353[19:0] ;
            mult_reg354[19:0] <= #DLY mult_wire354[19:0] ;
            mult_reg355[19:0] <= #DLY mult_wire355[19:0] ;
            mult_reg356[19:0] <= #DLY mult_wire356[19:0] ;
            mult_reg357[19:0] <= #DLY mult_wire357[19:0] ;
            mult_reg358[19:0] <= #DLY mult_wire358[19:0] ;
            mult_reg359[19:0] <= #DLY mult_wire359[19:0] ;
            mult_reg360[19:0] <= #DLY mult_wire360[19:0] ;
            mult_reg361[19:0] <= #DLY mult_wire361[19:0] ;
            mult_reg362[19:0] <= #DLY mult_wire362[19:0] ;
            mult_reg363[19:0] <= #DLY mult_wire363[19:0] ;
            mult_reg364[19:0] <= #DLY mult_wire364[19:0] ;
            mult_reg365[19:0] <= #DLY mult_wire365[19:0] ;
            mult_reg366[19:0] <= #DLY mult_wire366[19:0] ;
            mult_reg367[19:0] <= #DLY mult_wire367[19:0] ;
            mult_reg368[19:0] <= #DLY mult_wire368[19:0] ;
            mult_reg369[19:0] <= #DLY mult_wire369[19:0] ;
            mult_reg370[19:0] <= #DLY mult_wire370[19:0] ;
            mult_reg371[19:0] <= #DLY mult_wire371[19:0] ;
            mult_reg372[19:0] <= #DLY mult_wire372[19:0] ;
            mult_reg373[19:0] <= #DLY mult_wire373[19:0] ;
            mult_reg374[19:0] <= #DLY mult_wire374[19:0] ;
            mult_reg375[19:0] <= #DLY mult_wire375[19:0] ;
            mult_reg376[19:0] <= #DLY mult_wire376[19:0] ;
            mult_reg377[19:0] <= #DLY mult_wire377[19:0] ;
            mult_reg378[19:0] <= #DLY mult_wire378[19:0] ;
            mult_reg379[19:0] <= #DLY mult_wire379[19:0] ;
            mult_reg380[19:0] <= #DLY mult_wire380[19:0] ;
            mult_reg381[19:0] <= #DLY mult_wire381[19:0] ;
            mult_reg382[19:0] <= #DLY mult_wire382[19:0] ;
            mult_reg383[19:0] <= #DLY mult_wire383[19:0] ;
            mult_reg384[19:0] <= #DLY mult_wire384[19:0] ;
            mult_reg385[19:0] <= #DLY mult_wire385[19:0] ;
            mult_reg386[19:0] <= #DLY mult_wire386[19:0] ;
            mult_reg387[19:0] <= #DLY mult_wire387[19:0] ;
            mult_reg388[19:0] <= #DLY mult_wire388[19:0] ;
            mult_reg389[19:0] <= #DLY mult_wire389[19:0] ;
            mult_reg390[19:0] <= #DLY mult_wire390[19:0] ;
            mult_reg391[19:0] <= #DLY mult_wire391[19:0] ;
            mult_reg392[19:0] <= #DLY mult_wire392[19:0] ;
            mult_reg393[19:0] <= #DLY mult_wire393[19:0] ;
            mult_reg394[19:0] <= #DLY mult_wire394[19:0] ;
            mult_reg395[19:0] <= #DLY mult_wire395[19:0] ;
            mult_reg396[19:0] <= #DLY mult_wire396[19:0] ;
            mult_reg397[19:0] <= #DLY mult_wire397[19:0] ;
            mult_reg398[19:0] <= #DLY mult_wire398[19:0] ;
            mult_reg399[19:0] <= #DLY mult_wire399[19:0] ;
            mult_reg400[19:0] <= #DLY mult_wire400[19:0] ;
            mult_reg401[19:0] <= #DLY mult_wire401[19:0] ;
            mult_reg402[19:0] <= #DLY mult_wire402[19:0] ;
            mult_reg403[19:0] <= #DLY mult_wire403[19:0] ;
            mult_reg404[19:0] <= #DLY mult_wire404[19:0] ;
            mult_reg405[19:0] <= #DLY mult_wire405[19:0] ;
            mult_reg406[19:0] <= #DLY mult_wire406[19:0] ;
            mult_reg407[19:0] <= #DLY mult_wire407[19:0] ;
            mult_reg408[19:0] <= #DLY mult_wire408[19:0] ;
            mult_reg409[19:0] <= #DLY mult_wire409[19:0] ;
            mult_reg410[19:0] <= #DLY mult_wire410[19:0] ;
            mult_reg411[19:0] <= #DLY mult_wire411[19:0] ;
            mult_reg412[19:0] <= #DLY mult_wire412[19:0] ;
            mult_reg413[19:0] <= #DLY mult_wire413[19:0] ;
            mult_reg414[19:0] <= #DLY mult_wire414[19:0] ;
            mult_reg415[19:0] <= #DLY mult_wire415[19:0] ;
            mult_reg416[19:0] <= #DLY mult_wire416[19:0] ;
            mult_reg417[19:0] <= #DLY mult_wire417[19:0] ;
            mult_reg418[19:0] <= #DLY mult_wire418[19:0] ;
            mult_reg419[19:0] <= #DLY mult_wire419[19:0] ;
            mult_reg420[19:0] <= #DLY mult_wire420[19:0] ;
            mult_reg421[19:0] <= #DLY mult_wire421[19:0] ;
            mult_reg422[19:0] <= #DLY mult_wire422[19:0] ;
            mult_reg423[19:0] <= #DLY mult_wire423[19:0] ;
            mult_reg424[19:0] <= #DLY mult_wire424[19:0] ;
            mult_reg425[19:0] <= #DLY mult_wire425[19:0] ;
            mult_reg426[19:0] <= #DLY mult_wire426[19:0] ;
            mult_reg427[19:0] <= #DLY mult_wire427[19:0] ;
            mult_reg428[19:0] <= #DLY mult_wire428[19:0] ;
            mult_reg429[19:0] <= #DLY mult_wire429[19:0] ;
            mult_reg430[19:0] <= #DLY mult_wire430[19:0] ;
            mult_reg431[19:0] <= #DLY mult_wire431[19:0] ;
            mult_reg432[19:0] <= #DLY mult_wire432[19:0] ;
            mult_reg433[19:0] <= #DLY mult_wire433[19:0] ;
            mult_reg434[19:0] <= #DLY mult_wire434[19:0] ;
            mult_reg435[19:0] <= #DLY mult_wire435[19:0] ;
            mult_reg436[19:0] <= #DLY mult_wire436[19:0] ;
            mult_reg437[19:0] <= #DLY mult_wire437[19:0] ;
            mult_reg438[19:0] <= #DLY mult_wire438[19:0] ;
            mult_reg439[19:0] <= #DLY mult_wire439[19:0] ;
            mult_reg440[19:0] <= #DLY mult_wire440[19:0] ;
            mult_reg441[19:0] <= #DLY mult_wire441[19:0] ;
            mult_reg442[19:0] <= #DLY mult_wire442[19:0] ;
            mult_reg443[19:0] <= #DLY mult_wire443[19:0] ;
            mult_reg444[19:0] <= #DLY mult_wire444[19:0] ;
            mult_reg445[19:0] <= #DLY mult_wire445[19:0] ;
            mult_reg446[19:0] <= #DLY mult_wire446[19:0] ;
            mult_reg447[19:0] <= #DLY mult_wire447[19:0] ;
            mult_reg448[19:0] <= #DLY mult_wire448[19:0] ;
            mult_reg449[19:0] <= #DLY mult_wire449[19:0] ;
            mult_reg450[19:0] <= #DLY mult_wire450[19:0] ;
            mult_reg451[19:0] <= #DLY mult_wire451[19:0] ;
            mult_reg452[19:0] <= #DLY mult_wire452[19:0] ;
            mult_reg453[19:0] <= #DLY mult_wire453[19:0] ;
            mult_reg454[19:0] <= #DLY mult_wire454[19:0] ;
            mult_reg455[19:0] <= #DLY mult_wire455[19:0] ;
            mult_reg456[19:0] <= #DLY mult_wire456[19:0] ;
            mult_reg457[19:0] <= #DLY mult_wire457[19:0] ;
            mult_reg458[19:0] <= #DLY mult_wire458[19:0] ;
            mult_reg459[19:0] <= #DLY mult_wire459[19:0] ;
            mult_reg460[19:0] <= #DLY mult_wire460[19:0] ;
            mult_reg461[19:0] <= #DLY mult_wire461[19:0] ;
            mult_reg462[19:0] <= #DLY mult_wire462[19:0] ;
            mult_reg463[19:0] <= #DLY mult_wire463[19:0] ;
            mult_reg464[19:0] <= #DLY mult_wire464[19:0] ;
            mult_reg465[19:0] <= #DLY mult_wire465[19:0] ;
            mult_reg466[19:0] <= #DLY mult_wire466[19:0] ;
            mult_reg467[19:0] <= #DLY mult_wire467[19:0] ;
            mult_reg468[19:0] <= #DLY mult_wire468[19:0] ;
            mult_reg469[19:0] <= #DLY mult_wire469[19:0] ;
            mult_reg470[19:0] <= #DLY mult_wire470[19:0] ;
            mult_reg471[19:0] <= #DLY mult_wire471[19:0] ;
            mult_reg472[19:0] <= #DLY mult_wire472[19:0] ;
            mult_reg473[19:0] <= #DLY mult_wire473[19:0] ;
            mult_reg474[19:0] <= #DLY mult_wire474[19:0] ;
            mult_reg475[19:0] <= #DLY mult_wire475[19:0] ;
            mult_reg476[19:0] <= #DLY mult_wire476[19:0] ;
            mult_reg477[19:0] <= #DLY mult_wire477[19:0] ;
            mult_reg478[19:0] <= #DLY mult_wire478[19:0] ;
            mult_reg479[19:0] <= #DLY mult_wire479[19:0] ;
            mult_reg480[19:0] <= #DLY mult_wire480[19:0] ;
            mult_reg481[19:0] <= #DLY mult_wire481[19:0] ;
            mult_reg482[19:0] <= #DLY mult_wire482[19:0] ;
            mult_reg483[19:0] <= #DLY mult_wire483[19:0] ;
            mult_reg484[19:0] <= #DLY mult_wire484[19:0] ;
            mult_reg485[19:0] <= #DLY mult_wire485[19:0] ;
            mult_reg486[19:0] <= #DLY mult_wire486[19:0] ;
            mult_reg487[19:0] <= #DLY mult_wire487[19:0] ;
            mult_reg488[19:0] <= #DLY mult_wire488[19:0] ;
            mult_reg489[19:0] <= #DLY mult_wire489[19:0] ;
            mult_reg490[19:0] <= #DLY mult_wire490[19:0] ;
            mult_reg491[19:0] <= #DLY mult_wire491[19:0] ;
            mult_reg492[19:0] <= #DLY mult_wire492[19:0] ;
            mult_reg493[19:0] <= #DLY mult_wire493[19:0] ;
            mult_reg494[19:0] <= #DLY mult_wire494[19:0] ;
            mult_reg495[19:0] <= #DLY mult_wire495[19:0] ;
            mult_reg496[19:0] <= #DLY mult_wire496[19:0] ;
            mult_reg497[19:0] <= #DLY mult_wire497[19:0] ;
            mult_reg498[19:0] <= #DLY mult_wire498[19:0] ;
            mult_reg499[19:0] <= #DLY mult_wire499[19:0] ;
            mult_reg500[19:0] <= #DLY mult_wire500[19:0] ;
            mult_reg501[19:0] <= #DLY mult_wire501[19:0] ;
            mult_reg502[19:0] <= #DLY mult_wire502[19:0] ;
            mult_reg503[19:0] <= #DLY mult_wire503[19:0] ;
            mult_reg504[19:0] <= #DLY mult_wire504[19:0] ;
            mult_reg505[19:0] <= #DLY mult_wire505[19:0] ;
            mult_reg506[19:0] <= #DLY mult_wire506[19:0] ;
            mult_reg507[19:0] <= #DLY mult_wire507[19:0] ;
            mult_reg508[19:0] <= #DLY mult_wire508[19:0] ;
            mult_reg509[19:0] <= #DLY mult_wire509[19:0] ;
            mult_reg510[19:0] <= #DLY mult_wire510[19:0] ;
            mult_reg511[19:0] <= #DLY mult_wire511[19:0] ;
            mult_reg512[19:0] <= #DLY mult_wire512[19:0] ;
		end
	end

    /****************************
    // pipeline[34] Active
    ****************************/
    wire [20:0] sum512_256_wire01  = {1'd0, mult_reg01[19:0]}  + {1'd0, mult_reg02[19:0]}  ;
    wire [20:0] sum512_256_wire02  = {1'd0, mult_reg03[19:0]}  + {1'd0, mult_reg04[19:0]}  ;
    wire [20:0] sum512_256_wire03  = {1'd0, mult_reg05[19:0]}  + {1'd0, mult_reg06[19:0]}  ;
    wire [20:0] sum512_256_wire04  = {1'd0, mult_reg07[19:0]}  + {1'd0, mult_reg08[19:0]}  ;
    wire [20:0] sum512_256_wire05  = {1'd0, mult_reg09[19:0]}  + {1'd0, mult_reg10[19:0]}  ;
    wire [20:0] sum512_256_wire06  = {1'd0, mult_reg11[19:0]}  + {1'd0, mult_reg12[19:0]}  ;
    wire [20:0] sum512_256_wire07  = {1'd0, mult_reg13[19:0]}  + {1'd0, mult_reg14[19:0]}  ;
    wire [20:0] sum512_256_wire08  = {1'd0, mult_reg15[19:0]}  + {1'd0, mult_reg16[19:0]}  ;
    wire [20:0] sum512_256_wire09  = {1'd0, mult_reg17[19:0]}  + {1'd0, mult_reg18[19:0]}  ;
    wire [20:0] sum512_256_wire10  = {1'd0, mult_reg19[19:0]}  + {1'd0, mult_reg20[19:0]}  ;
    wire [20:0] sum512_256_wire11  = {1'd0, mult_reg21[19:0]}  + {1'd0, mult_reg22[19:0]}  ;
    wire [20:0] sum512_256_wire12  = {1'd0, mult_reg23[19:0]}  + {1'd0, mult_reg24[19:0]}  ;
    wire [20:0] sum512_256_wire13  = {1'd0, mult_reg25[19:0]}  + {1'd0, mult_reg26[19:0]}  ;
    wire [20:0] sum512_256_wire14  = {1'd0, mult_reg27[19:0]}  + {1'd0, mult_reg28[19:0]}  ;
    wire [20:0] sum512_256_wire15  = {1'd0, mult_reg29[19:0]}  + {1'd0, mult_reg30[19:0]}  ;
    wire [20:0] sum512_256_wire16  = {1'd0, mult_reg31[19:0]}  + {1'd0, mult_reg32[19:0]}  ;
    wire [20:0] sum512_256_wire17  = {1'd0, mult_reg33[19:0]}  + {1'd0, mult_reg34[19:0]}  ;
    wire [20:0] sum512_256_wire18  = {1'd0, mult_reg35[19:0]}  + {1'd0, mult_reg36[19:0]}  ;
    wire [20:0] sum512_256_wire19  = {1'd0, mult_reg37[19:0]}  + {1'd0, mult_reg38[19:0]}  ;
    wire [20:0] sum512_256_wire20  = {1'd0, mult_reg39[19:0]}  + {1'd0, mult_reg40[19:0]}  ;
    wire [20:0] sum512_256_wire21  = {1'd0, mult_reg41[19:0]}  + {1'd0, mult_reg42[19:0]}  ;
    wire [20:0] sum512_256_wire22  = {1'd0, mult_reg43[19:0]}  + {1'd0, mult_reg44[19:0]}  ;
    wire [20:0] sum512_256_wire23  = {1'd0, mult_reg45[19:0]}  + {1'd0, mult_reg46[19:0]}  ;
    wire [20:0] sum512_256_wire24  = {1'd0, mult_reg47[19:0]}  + {1'd0, mult_reg48[19:0]}  ;
    wire [20:0] sum512_256_wire25  = {1'd0, mult_reg49[19:0]}  + {1'd0, mult_reg50[19:0]}  ;
    wire [20:0] sum512_256_wire26  = {1'd0, mult_reg51[19:0]}  + {1'd0, mult_reg52[19:0]}  ;
    wire [20:0] sum512_256_wire27  = {1'd0, mult_reg53[19:0]}  + {1'd0, mult_reg54[19:0]}  ;
    wire [20:0] sum512_256_wire28  = {1'd0, mult_reg55[19:0]}  + {1'd0, mult_reg56[19:0]}  ;
    wire [20:0] sum512_256_wire29  = {1'd0, mult_reg57[19:0]}  + {1'd0, mult_reg58[19:0]}  ;
    wire [20:0] sum512_256_wire30  = {1'd0, mult_reg59[19:0]}  + {1'd0, mult_reg60[19:0]}  ;
    wire [20:0] sum512_256_wire31  = {1'd0, mult_reg61[19:0]}  + {1'd0, mult_reg62[19:0]}  ;
    wire [20:0] sum512_256_wire32  = {1'd0, mult_reg63[19:0]}  + {1'd0, mult_reg64[19:0]}  ;
    wire [20:0] sum512_256_wire33  = {1'd0, mult_reg65[19:0]}  + {1'd0, mult_reg66[19:0]}  ;
    wire [20:0] sum512_256_wire34  = {1'd0, mult_reg67[19:0]}  + {1'd0, mult_reg68[19:0]}  ;
    wire [20:0] sum512_256_wire35  = {1'd0, mult_reg69[19:0]}  + {1'd0, mult_reg70[19:0]}  ;
    wire [20:0] sum512_256_wire36  = {1'd0, mult_reg71[19:0]}  + {1'd0, mult_reg72[19:0]}  ;
    wire [20:0] sum512_256_wire37  = {1'd0, mult_reg73[19:0]}  + {1'd0, mult_reg74[19:0]}  ;
    wire [20:0] sum512_256_wire38  = {1'd0, mult_reg75[19:0]}  + {1'd0, mult_reg76[19:0]}  ;
    wire [20:0] sum512_256_wire39  = {1'd0, mult_reg77[19:0]}  + {1'd0, mult_reg78[19:0]}  ;
    wire [20:0] sum512_256_wire40  = {1'd0, mult_reg79[19:0]}  + {1'd0, mult_reg80[19:0]}  ;
    wire [20:0] sum512_256_wire41  = {1'd0, mult_reg81[19:0]}  + {1'd0, mult_reg82[19:0]}  ;
    wire [20:0] sum512_256_wire42  = {1'd0, mult_reg83[19:0]}  + {1'd0, mult_reg84[19:0]}  ;
    wire [20:0] sum512_256_wire43  = {1'd0, mult_reg85[19:0]}  + {1'd0, mult_reg86[19:0]}  ;
    wire [20:0] sum512_256_wire44  = {1'd0, mult_reg87[19:0]}  + {1'd0, mult_reg88[19:0]}  ;
    wire [20:0] sum512_256_wire45  = {1'd0, mult_reg89[19:0]}  + {1'd0, mult_reg90[19:0]}  ;
    wire [20:0] sum512_256_wire46  = {1'd0, mult_reg91[19:0]}  + {1'd0, mult_reg92[19:0]}  ;
    wire [20:0] sum512_256_wire47  = {1'd0, mult_reg93[19:0]}  + {1'd0, mult_reg94[19:0]}  ;
    wire [20:0] sum512_256_wire48  = {1'd0, mult_reg95[19:0]}  + {1'd0, mult_reg96[19:0]}  ;
    wire [20:0] sum512_256_wire49  = {1'd0, mult_reg97[19:0]}  + {1'd0, mult_reg98[19:0]}  ;
    wire [20:0] sum512_256_wire50  = {1'd0, mult_reg99[19:0]}  + {1'd0, mult_reg100[19:0]} ;
    wire [20:0] sum512_256_wire51  = {1'd0, mult_reg101[19:0]} + {1'd0, mult_reg102[19:0]} ;
    wire [20:0] sum512_256_wire52  = {1'd0, mult_reg103[19:0]} + {1'd0, mult_reg104[19:0]} ;
    wire [20:0] sum512_256_wire53  = {1'd0, mult_reg105[19:0]} + {1'd0, mult_reg106[19:0]} ;
    wire [20:0] sum512_256_wire54  = {1'd0, mult_reg107[19:0]} + {1'd0, mult_reg108[19:0]} ;
    wire [20:0] sum512_256_wire55  = {1'd0, mult_reg109[19:0]} + {1'd0, mult_reg110[19:0]} ;
    wire [20:0] sum512_256_wire56  = {1'd0, mult_reg111[19:0]} + {1'd0, mult_reg112[19:0]} ;
    wire [20:0] sum512_256_wire57  = {1'd0, mult_reg113[19:0]} + {1'd0, mult_reg114[19:0]} ;
    wire [20:0] sum512_256_wire58  = {1'd0, mult_reg115[19:0]} + {1'd0, mult_reg116[19:0]} ;
    wire [20:0] sum512_256_wire59  = {1'd0, mult_reg117[19:0]} + {1'd0, mult_reg118[19:0]} ;
    wire [20:0] sum512_256_wire60  = {1'd0, mult_reg119[19:0]} + {1'd0, mult_reg120[19:0]} ;
    wire [20:0] sum512_256_wire61  = {1'd0, mult_reg121[19:0]} + {1'd0, mult_reg122[19:0]} ;
    wire [20:0] sum512_256_wire62  = {1'd0, mult_reg123[19:0]} + {1'd0, mult_reg124[19:0]} ;
    wire [20:0] sum512_256_wire63  = {1'd0, mult_reg125[19:0]} + {1'd0, mult_reg126[19:0]} ;
    wire [20:0] sum512_256_wire64  = {1'd0, mult_reg127[19:0]} + {1'd0, mult_reg128[19:0]} ;
    wire [20:0] sum512_256_wire65  = {1'd0, mult_reg129[19:0]} + {1'd0, mult_reg130[19:0]} ;
    wire [20:0] sum512_256_wire66  = {1'd0, mult_reg131[19:0]} + {1'd0, mult_reg132[19:0]} ;
    wire [20:0] sum512_256_wire67  = {1'd0, mult_reg133[19:0]} + {1'd0, mult_reg134[19:0]} ;
    wire [20:0] sum512_256_wire68  = {1'd0, mult_reg135[19:0]} + {1'd0, mult_reg136[19:0]} ;
    wire [20:0] sum512_256_wire69  = {1'd0, mult_reg137[19:0]} + {1'd0, mult_reg138[19:0]} ;
    wire [20:0] sum512_256_wire70  = {1'd0, mult_reg139[19:0]} + {1'd0, mult_reg140[19:0]} ;
    wire [20:0] sum512_256_wire71  = {1'd0, mult_reg141[19:0]} + {1'd0, mult_reg142[19:0]} ;
    wire [20:0] sum512_256_wire72  = {1'd0, mult_reg143[19:0]} + {1'd0, mult_reg144[19:0]} ;
    wire [20:0] sum512_256_wire73  = {1'd0, mult_reg145[19:0]} + {1'd0, mult_reg146[19:0]} ;
    wire [20:0] sum512_256_wire74  = {1'd0, mult_reg147[19:0]} + {1'd0, mult_reg148[19:0]} ;
    wire [20:0] sum512_256_wire75  = {1'd0, mult_reg149[19:0]} + {1'd0, mult_reg150[19:0]} ;
    wire [20:0] sum512_256_wire76  = {1'd0, mult_reg151[19:0]} + {1'd0, mult_reg152[19:0]} ;
    wire [20:0] sum512_256_wire77  = {1'd0, mult_reg153[19:0]} + {1'd0, mult_reg154[19:0]} ;
    wire [20:0] sum512_256_wire78  = {1'd0, mult_reg155[19:0]} + {1'd0, mult_reg156[19:0]} ;
    wire [20:0] sum512_256_wire79  = {1'd0, mult_reg157[19:0]} + {1'd0, mult_reg158[19:0]} ;
    wire [20:0] sum512_256_wire80  = {1'd0, mult_reg159[19:0]} + {1'd0, mult_reg160[19:0]} ;
    wire [20:0] sum512_256_wire81  = {1'd0, mult_reg161[19:0]} + {1'd0, mult_reg162[19:0]} ;
    wire [20:0] sum512_256_wire82  = {1'd0, mult_reg163[19:0]} + {1'd0, mult_reg164[19:0]} ;
    wire [20:0] sum512_256_wire83  = {1'd0, mult_reg165[19:0]} + {1'd0, mult_reg166[19:0]} ;
    wire [20:0] sum512_256_wire84  = {1'd0, mult_reg167[19:0]} + {1'd0, mult_reg168[19:0]} ;
    wire [20:0] sum512_256_wire85  = {1'd0, mult_reg169[19:0]} + {1'd0, mult_reg170[19:0]} ;
    wire [20:0] sum512_256_wire86  = {1'd0, mult_reg171[19:0]} + {1'd0, mult_reg172[19:0]} ;
    wire [20:0] sum512_256_wire87  = {1'd0, mult_reg173[19:0]} + {1'd0, mult_reg174[19:0]} ;
    wire [20:0] sum512_256_wire88  = {1'd0, mult_reg175[19:0]} + {1'd0, mult_reg176[19:0]} ;
    wire [20:0] sum512_256_wire89  = {1'd0, mult_reg177[19:0]} + {1'd0, mult_reg178[19:0]} ;
    wire [20:0] sum512_256_wire90  = {1'd0, mult_reg179[19:0]} + {1'd0, mult_reg180[19:0]} ;
    wire [20:0] sum512_256_wire91  = {1'd0, mult_reg181[19:0]} + {1'd0, mult_reg182[19:0]} ;
    wire [20:0] sum512_256_wire92  = {1'd0, mult_reg183[19:0]} + {1'd0, mult_reg184[19:0]} ;
    wire [20:0] sum512_256_wire93  = {1'd0, mult_reg185[19:0]} + {1'd0, mult_reg186[19:0]} ;
    wire [20:0] sum512_256_wire94  = {1'd0, mult_reg187[19:0]} + {1'd0, mult_reg188[19:0]} ;
    wire [20:0] sum512_256_wire95  = {1'd0, mult_reg189[19:0]} + {1'd0, mult_reg190[19:0]} ;
    wire [20:0] sum512_256_wire96  = {1'd0, mult_reg191[19:0]} + {1'd0, mult_reg192[19:0]} ;
    wire [20:0] sum512_256_wire97  = {1'd0, mult_reg193[19:0]} + {1'd0, mult_reg194[19:0]} ;
    wire [20:0] sum512_256_wire98  = {1'd0, mult_reg195[19:0]} + {1'd0, mult_reg196[19:0]} ;
    wire [20:0] sum512_256_wire99  = {1'd0, mult_reg197[19:0]} + {1'd0, mult_reg198[19:0]} ;
    wire [20:0] sum512_256_wire100 = {1'd0, mult_reg199[19:0]} + {1'd0, mult_reg200[19:0]} ;
    wire [20:0] sum512_256_wire101 = {1'd0, mult_reg201[19:0]} + {1'd0, mult_reg202[19:0]} ;
    wire [20:0] sum512_256_wire102 = {1'd0, mult_reg203[19:0]} + {1'd0, mult_reg204[19:0]} ;
    wire [20:0] sum512_256_wire103 = {1'd0, mult_reg205[19:0]} + {1'd0, mult_reg206[19:0]} ;
    wire [20:0] sum512_256_wire104 = {1'd0, mult_reg207[19:0]} + {1'd0, mult_reg208[19:0]} ;
    wire [20:0] sum512_256_wire105 = {1'd0, mult_reg209[19:0]} + {1'd0, mult_reg210[19:0]} ;
    wire [20:0] sum512_256_wire106 = {1'd0, mult_reg211[19:0]} + {1'd0, mult_reg212[19:0]} ;
    wire [20:0] sum512_256_wire107 = {1'd0, mult_reg213[19:0]} + {1'd0, mult_reg214[19:0]} ;
    wire [20:0] sum512_256_wire108 = {1'd0, mult_reg215[19:0]} + {1'd0, mult_reg216[19:0]} ;
    wire [20:0] sum512_256_wire109 = {1'd0, mult_reg217[19:0]} + {1'd0, mult_reg218[19:0]} ;
    wire [20:0] sum512_256_wire110 = {1'd0, mult_reg219[19:0]} + {1'd0, mult_reg220[19:0]} ;
    wire [20:0] sum512_256_wire111 = {1'd0, mult_reg221[19:0]} + {1'd0, mult_reg222[19:0]} ;
    wire [20:0] sum512_256_wire112 = {1'd0, mult_reg223[19:0]} + {1'd0, mult_reg224[19:0]} ;
    wire [20:0] sum512_256_wire113 = {1'd0, mult_reg225[19:0]} + {1'd0, mult_reg226[19:0]} ;
    wire [20:0] sum512_256_wire114 = {1'd0, mult_reg227[19:0]} + {1'd0, mult_reg228[19:0]} ;
    wire [20:0] sum512_256_wire115 = {1'd0, mult_reg229[19:0]} + {1'd0, mult_reg230[19:0]} ;
    wire [20:0] sum512_256_wire116 = {1'd0, mult_reg231[19:0]} + {1'd0, mult_reg232[19:0]} ;
    wire [20:0] sum512_256_wire117 = {1'd0, mult_reg233[19:0]} + {1'd0, mult_reg234[19:0]} ;
    wire [20:0] sum512_256_wire118 = {1'd0, mult_reg235[19:0]} + {1'd0, mult_reg236[19:0]} ;
    wire [20:0] sum512_256_wire119 = {1'd0, mult_reg237[19:0]} + {1'd0, mult_reg238[19:0]} ;
    wire [20:0] sum512_256_wire120 = {1'd0, mult_reg239[19:0]} + {1'd0, mult_reg240[19:0]} ;
    wire [20:0] sum512_256_wire121 = {1'd0, mult_reg241[19:0]} + {1'd0, mult_reg242[19:0]} ;
    wire [20:0] sum512_256_wire122 = {1'd0, mult_reg243[19:0]} + {1'd0, mult_reg244[19:0]} ;
    wire [20:0] sum512_256_wire123 = {1'd0, mult_reg245[19:0]} + {1'd0, mult_reg246[19:0]} ;
    wire [20:0] sum512_256_wire124 = {1'd0, mult_reg247[19:0]} + {1'd0, mult_reg248[19:0]} ;
    wire [20:0] sum512_256_wire125 = {1'd0, mult_reg249[19:0]} + {1'd0, mult_reg250[19:0]} ;
    wire [20:0] sum512_256_wire126 = {1'd0, mult_reg251[19:0]} + {1'd0, mult_reg252[19:0]} ;
    wire [20:0] sum512_256_wire127 = {1'd0, mult_reg253[19:0]} + {1'd0, mult_reg254[19:0]} ;
    wire [20:0] sum512_256_wire128 = {1'd0, mult_reg255[19:0]} + {1'd0, mult_reg256[19:0]} ;
    wire [20:0] sum512_256_wire129 = {1'd0, mult_reg257[19:0]} + {1'd0, mult_reg258[19:0]} ;
    wire [20:0] sum512_256_wire130 = {1'd0, mult_reg259[19:0]} + {1'd0, mult_reg260[19:0]} ;
    wire [20:0] sum512_256_wire131 = {1'd0, mult_reg261[19:0]} + {1'd0, mult_reg262[19:0]} ;
    wire [20:0] sum512_256_wire132 = {1'd0, mult_reg263[19:0]} + {1'd0, mult_reg264[19:0]} ;
    wire [20:0] sum512_256_wire133 = {1'd0, mult_reg265[19:0]} + {1'd0, mult_reg266[19:0]} ;
    wire [20:0] sum512_256_wire134 = {1'd0, mult_reg267[19:0]} + {1'd0, mult_reg268[19:0]} ;
    wire [20:0] sum512_256_wire135 = {1'd0, mult_reg269[19:0]} + {1'd0, mult_reg270[19:0]} ;
    wire [20:0] sum512_256_wire136 = {1'd0, mult_reg271[19:0]} + {1'd0, mult_reg272[19:0]} ;
    wire [20:0] sum512_256_wire137 = {1'd0, mult_reg273[19:0]} + {1'd0, mult_reg274[19:0]} ;
    wire [20:0] sum512_256_wire138 = {1'd0, mult_reg275[19:0]} + {1'd0, mult_reg276[19:0]} ;
    wire [20:0] sum512_256_wire139 = {1'd0, mult_reg277[19:0]} + {1'd0, mult_reg278[19:0]} ;
    wire [20:0] sum512_256_wire140 = {1'd0, mult_reg279[19:0]} + {1'd0, mult_reg280[19:0]} ;
    wire [20:0] sum512_256_wire141 = {1'd0, mult_reg281[19:0]} + {1'd0, mult_reg282[19:0]} ;
    wire [20:0] sum512_256_wire142 = {1'd0, mult_reg283[19:0]} + {1'd0, mult_reg284[19:0]} ;
    wire [20:0] sum512_256_wire143 = {1'd0, mult_reg285[19:0]} + {1'd0, mult_reg286[19:0]} ;
    wire [20:0] sum512_256_wire144 = {1'd0, mult_reg287[19:0]} + {1'd0, mult_reg288[19:0]} ;
    wire [20:0] sum512_256_wire145 = {1'd0, mult_reg289[19:0]} + {1'd0, mult_reg290[19:0]} ;
    wire [20:0] sum512_256_wire146 = {1'd0, mult_reg291[19:0]} + {1'd0, mult_reg292[19:0]} ;
    wire [20:0] sum512_256_wire147 = {1'd0, mult_reg293[19:0]} + {1'd0, mult_reg294[19:0]} ;
    wire [20:0] sum512_256_wire148 = {1'd0, mult_reg295[19:0]} + {1'd0, mult_reg296[19:0]} ;
    wire [20:0] sum512_256_wire149 = {1'd0, mult_reg297[19:0]} + {1'd0, mult_reg298[19:0]} ;
    wire [20:0] sum512_256_wire150 = {1'd0, mult_reg299[19:0]} + {1'd0, mult_reg300[19:0]} ;
    wire [20:0] sum512_256_wire151 = {1'd0, mult_reg301[19:0]} + {1'd0, mult_reg302[19:0]} ;
    wire [20:0] sum512_256_wire152 = {1'd0, mult_reg303[19:0]} + {1'd0, mult_reg304[19:0]} ;
    wire [20:0] sum512_256_wire153 = {1'd0, mult_reg305[19:0]} + {1'd0, mult_reg306[19:0]} ;
    wire [20:0] sum512_256_wire154 = {1'd0, mult_reg307[19:0]} + {1'd0, mult_reg308[19:0]} ;
    wire [20:0] sum512_256_wire155 = {1'd0, mult_reg309[19:0]} + {1'd0, mult_reg310[19:0]} ;
    wire [20:0] sum512_256_wire156 = {1'd0, mult_reg311[19:0]} + {1'd0, mult_reg312[19:0]} ;
    wire [20:0] sum512_256_wire157 = {1'd0, mult_reg313[19:0]} + {1'd0, mult_reg314[19:0]} ;
    wire [20:0] sum512_256_wire158 = {1'd0, mult_reg315[19:0]} + {1'd0, mult_reg316[19:0]} ;
    wire [20:0] sum512_256_wire159 = {1'd0, mult_reg317[19:0]} + {1'd0, mult_reg318[19:0]} ;
    wire [20:0] sum512_256_wire160 = {1'd0, mult_reg319[19:0]} + {1'd0, mult_reg320[19:0]} ;
    wire [20:0] sum512_256_wire161 = {1'd0, mult_reg321[19:0]} + {1'd0, mult_reg322[19:0]} ;
    wire [20:0] sum512_256_wire162 = {1'd0, mult_reg323[19:0]} + {1'd0, mult_reg324[19:0]} ;
    wire [20:0] sum512_256_wire163 = {1'd0, mult_reg325[19:0]} + {1'd0, mult_reg326[19:0]} ;
    wire [20:0] sum512_256_wire164 = {1'd0, mult_reg327[19:0]} + {1'd0, mult_reg328[19:0]} ;
    wire [20:0] sum512_256_wire165 = {1'd0, mult_reg329[19:0]} + {1'd0, mult_reg330[19:0]} ;
    wire [20:0] sum512_256_wire166 = {1'd0, mult_reg331[19:0]} + {1'd0, mult_reg332[19:0]} ;
    wire [20:0] sum512_256_wire167 = {1'd0, mult_reg333[19:0]} + {1'd0, mult_reg334[19:0]} ;
    wire [20:0] sum512_256_wire168 = {1'd0, mult_reg335[19:0]} + {1'd0, mult_reg336[19:0]} ;
    wire [20:0] sum512_256_wire169 = {1'd0, mult_reg337[19:0]} + {1'd0, mult_reg338[19:0]} ;
    wire [20:0] sum512_256_wire170 = {1'd0, mult_reg339[19:0]} + {1'd0, mult_reg340[19:0]} ;
    wire [20:0] sum512_256_wire171 = {1'd0, mult_reg341[19:0]} + {1'd0, mult_reg342[19:0]} ;
    wire [20:0] sum512_256_wire172 = {1'd0, mult_reg343[19:0]} + {1'd0, mult_reg344[19:0]} ;
    wire [20:0] sum512_256_wire173 = {1'd0, mult_reg345[19:0]} + {1'd0, mult_reg346[19:0]} ;
    wire [20:0] sum512_256_wire174 = {1'd0, mult_reg347[19:0]} + {1'd0, mult_reg348[19:0]} ;
    wire [20:0] sum512_256_wire175 = {1'd0, mult_reg349[19:0]} + {1'd0, mult_reg350[19:0]} ;
    wire [20:0] sum512_256_wire176 = {1'd0, mult_reg351[19:0]} + {1'd0, mult_reg352[19:0]} ;
    wire [20:0] sum512_256_wire177 = {1'd0, mult_reg353[19:0]} + {1'd0, mult_reg354[19:0]} ;
    wire [20:0] sum512_256_wire178 = {1'd0, mult_reg355[19:0]} + {1'd0, mult_reg356[19:0]} ;
    wire [20:0] sum512_256_wire179 = {1'd0, mult_reg357[19:0]} + {1'd0, mult_reg358[19:0]} ;
    wire [20:0] sum512_256_wire180 = {1'd0, mult_reg359[19:0]} + {1'd0, mult_reg360[19:0]} ;
    wire [20:0] sum512_256_wire181 = {1'd0, mult_reg361[19:0]} + {1'd0, mult_reg362[19:0]} ;
    wire [20:0] sum512_256_wire182 = {1'd0, mult_reg363[19:0]} + {1'd0, mult_reg364[19:0]} ;
    wire [20:0] sum512_256_wire183 = {1'd0, mult_reg365[19:0]} + {1'd0, mult_reg366[19:0]} ;
    wire [20:0] sum512_256_wire184 = {1'd0, mult_reg367[19:0]} + {1'd0, mult_reg368[19:0]} ;
    wire [20:0] sum512_256_wire185 = {1'd0, mult_reg369[19:0]} + {1'd0, mult_reg370[19:0]} ;
    wire [20:0] sum512_256_wire186 = {1'd0, mult_reg371[19:0]} + {1'd0, mult_reg372[19:0]} ;
    wire [20:0] sum512_256_wire187 = {1'd0, mult_reg373[19:0]} + {1'd0, mult_reg374[19:0]} ;
    wire [20:0] sum512_256_wire188 = {1'd0, mult_reg375[19:0]} + {1'd0, mult_reg376[19:0]} ;
    wire [20:0] sum512_256_wire189 = {1'd0, mult_reg377[19:0]} + {1'd0, mult_reg378[19:0]} ;
    wire [20:0] sum512_256_wire190 = {1'd0, mult_reg379[19:0]} + {1'd0, mult_reg380[19:0]} ;
    wire [20:0] sum512_256_wire191 = {1'd0, mult_reg381[19:0]} + {1'd0, mult_reg382[19:0]} ;
    wire [20:0] sum512_256_wire192 = {1'd0, mult_reg383[19:0]} + {1'd0, mult_reg384[19:0]} ;
    wire [20:0] sum512_256_wire193 = {1'd0, mult_reg385[19:0]} + {1'd0, mult_reg386[19:0]} ;
    wire [20:0] sum512_256_wire194 = {1'd0, mult_reg387[19:0]} + {1'd0, mult_reg388[19:0]} ;
    wire [20:0] sum512_256_wire195 = {1'd0, mult_reg389[19:0]} + {1'd0, mult_reg390[19:0]} ;
    wire [20:0] sum512_256_wire196 = {1'd0, mult_reg391[19:0]} + {1'd0, mult_reg392[19:0]} ;
    wire [20:0] sum512_256_wire197 = {1'd0, mult_reg393[19:0]} + {1'd0, mult_reg394[19:0]} ;
    wire [20:0] sum512_256_wire198 = {1'd0, mult_reg395[19:0]} + {1'd0, mult_reg396[19:0]} ;
    wire [20:0] sum512_256_wire199 = {1'd0, mult_reg397[19:0]} + {1'd0, mult_reg398[19:0]} ;
    wire [20:0] sum512_256_wire200 = {1'd0, mult_reg399[19:0]} + {1'd0, mult_reg400[19:0]} ;
    wire [20:0] sum512_256_wire201 = {1'd0, mult_reg401[19:0]} + {1'd0, mult_reg402[19:0]} ;
    wire [20:0] sum512_256_wire202 = {1'd0, mult_reg403[19:0]} + {1'd0, mult_reg404[19:0]} ;
    wire [20:0] sum512_256_wire203 = {1'd0, mult_reg405[19:0]} + {1'd0, mult_reg406[19:0]} ;
    wire [20:0] sum512_256_wire204 = {1'd0, mult_reg407[19:0]} + {1'd0, mult_reg408[19:0]} ;
    wire [20:0] sum512_256_wire205 = {1'd0, mult_reg409[19:0]} + {1'd0, mult_reg410[19:0]} ;
    wire [20:0] sum512_256_wire206 = {1'd0, mult_reg411[19:0]} + {1'd0, mult_reg412[19:0]} ;
    wire [20:0] sum512_256_wire207 = {1'd0, mult_reg413[19:0]} + {1'd0, mult_reg414[19:0]} ;
    wire [20:0] sum512_256_wire208 = {1'd0, mult_reg415[19:0]} + {1'd0, mult_reg416[19:0]} ;
    wire [20:0] sum512_256_wire209 = {1'd0, mult_reg417[19:0]} + {1'd0, mult_reg418[19:0]} ;
    wire [20:0] sum512_256_wire210 = {1'd0, mult_reg419[19:0]} + {1'd0, mult_reg420[19:0]} ;
    wire [20:0] sum512_256_wire211 = {1'd0, mult_reg421[19:0]} + {1'd0, mult_reg422[19:0]} ;
    wire [20:0] sum512_256_wire212 = {1'd0, mult_reg423[19:0]} + {1'd0, mult_reg424[19:0]} ;
    wire [20:0] sum512_256_wire213 = {1'd0, mult_reg425[19:0]} + {1'd0, mult_reg426[19:0]} ;
    wire [20:0] sum512_256_wire214 = {1'd0, mult_reg427[19:0]} + {1'd0, mult_reg428[19:0]} ;
    wire [20:0] sum512_256_wire215 = {1'd0, mult_reg429[19:0]} + {1'd0, mult_reg430[19:0]} ;
    wire [20:0] sum512_256_wire216 = {1'd0, mult_reg431[19:0]} + {1'd0, mult_reg432[19:0]} ;
    wire [20:0] sum512_256_wire217 = {1'd0, mult_reg433[19:0]} + {1'd0, mult_reg434[19:0]} ;
    wire [20:0] sum512_256_wire218 = {1'd0, mult_reg435[19:0]} + {1'd0, mult_reg436[19:0]} ;
    wire [20:0] sum512_256_wire219 = {1'd0, mult_reg437[19:0]} + {1'd0, mult_reg438[19:0]} ;
    wire [20:0] sum512_256_wire220 = {1'd0, mult_reg439[19:0]} + {1'd0, mult_reg440[19:0]} ;
    wire [20:0] sum512_256_wire221 = {1'd0, mult_reg441[19:0]} + {1'd0, mult_reg442[19:0]} ;
    wire [20:0] sum512_256_wire222 = {1'd0, mult_reg443[19:0]} + {1'd0, mult_reg444[19:0]} ;
    wire [20:0] sum512_256_wire223 = {1'd0, mult_reg445[19:0]} + {1'd0, mult_reg446[19:0]} ;
    wire [20:0] sum512_256_wire224 = {1'd0, mult_reg447[19:0]} + {1'd0, mult_reg448[19:0]} ;
    wire [20:0] sum512_256_wire225 = {1'd0, mult_reg449[19:0]} + {1'd0, mult_reg450[19:0]} ;
    wire [20:0] sum512_256_wire226 = {1'd0, mult_reg451[19:0]} + {1'd0, mult_reg452[19:0]} ;
    wire [20:0] sum512_256_wire227 = {1'd0, mult_reg453[19:0]} + {1'd0, mult_reg454[19:0]} ;
    wire [20:0] sum512_256_wire228 = {1'd0, mult_reg455[19:0]} + {1'd0, mult_reg456[19:0]} ;
    wire [20:0] sum512_256_wire229 = {1'd0, mult_reg457[19:0]} + {1'd0, mult_reg458[19:0]} ;
    wire [20:0] sum512_256_wire230 = {1'd0, mult_reg459[19:0]} + {1'd0, mult_reg460[19:0]} ;
    wire [20:0] sum512_256_wire231 = {1'd0, mult_reg461[19:0]} + {1'd0, mult_reg462[19:0]} ;
    wire [20:0] sum512_256_wire232 = {1'd0, mult_reg463[19:0]} + {1'd0, mult_reg464[19:0]} ;
    wire [20:0] sum512_256_wire233 = {1'd0, mult_reg465[19:0]} + {1'd0, mult_reg466[19:0]} ;
    wire [20:0] sum512_256_wire234 = {1'd0, mult_reg467[19:0]} + {1'd0, mult_reg468[19:0]} ;
    wire [20:0] sum512_256_wire235 = {1'd0, mult_reg469[19:0]} + {1'd0, mult_reg470[19:0]} ;
    wire [20:0] sum512_256_wire236 = {1'd0, mult_reg471[19:0]} + {1'd0, mult_reg472[19:0]} ;
    wire [20:0] sum512_256_wire237 = {1'd0, mult_reg473[19:0]} + {1'd0, mult_reg474[19:0]} ;
    wire [20:0] sum512_256_wire238 = {1'd0, mult_reg475[19:0]} + {1'd0, mult_reg476[19:0]} ;
    wire [20:0] sum512_256_wire239 = {1'd0, mult_reg477[19:0]} + {1'd0, mult_reg478[19:0]} ;
    wire [20:0] sum512_256_wire240 = {1'd0, mult_reg479[19:0]} + {1'd0, mult_reg480[19:0]} ;
    wire [20:0] sum512_256_wire241 = {1'd0, mult_reg481[19:0]} + {1'd0, mult_reg482[19:0]} ;
    wire [20:0] sum512_256_wire242 = {1'd0, mult_reg483[19:0]} + {1'd0, mult_reg484[19:0]} ;
    wire [20:0] sum512_256_wire243 = {1'd0, mult_reg485[19:0]} + {1'd0, mult_reg486[19:0]} ;
    wire [20:0] sum512_256_wire244 = {1'd0, mult_reg487[19:0]} + {1'd0, mult_reg488[19:0]} ;
    wire [20:0] sum512_256_wire245 = {1'd0, mult_reg489[19:0]} + {1'd0, mult_reg490[19:0]} ;
    wire [20:0] sum512_256_wire246 = {1'd0, mult_reg491[19:0]} + {1'd0, mult_reg492[19:0]} ;
    wire [20:0] sum512_256_wire247 = {1'd0, mult_reg493[19:0]} + {1'd0, mult_reg494[19:0]} ;
    wire [20:0] sum512_256_wire248 = {1'd0, mult_reg495[19:0]} + {1'd0, mult_reg496[19:0]} ;
    wire [20:0] sum512_256_wire249 = {1'd0, mult_reg497[19:0]} + {1'd0, mult_reg498[19:0]} ;
    wire [20:0] sum512_256_wire250 = {1'd0, mult_reg499[19:0]} + {1'd0, mult_reg500[19:0]} ;
    wire [20:0] sum512_256_wire251 = {1'd0, mult_reg501[19:0]} + {1'd0, mult_reg502[19:0]} ;
    wire [20:0] sum512_256_wire252 = {1'd0, mult_reg503[19:0]} + {1'd0, mult_reg504[19:0]} ;
    wire [20:0] sum512_256_wire253 = {1'd0, mult_reg505[19:0]} + {1'd0, mult_reg506[19:0]} ;
    wire [20:0] sum512_256_wire254 = {1'd0, mult_reg507[19:0]} + {1'd0, mult_reg508[19:0]} ;
    wire [20:0] sum512_256_wire255 = {1'd0, mult_reg509[19:0]} + {1'd0, mult_reg510[19:0]} ;
    wire [20:0] sum512_256_wire256 = {1'd0, mult_reg511[19:0]} + {1'd0, mult_reg512[19:0]} ;
    
    wire [21:0] sum256_128_wire01  = {1'd0, sum512_256_wire01[20:0]}  + {1'd0, sum512_256_wire02[20:0]}  ;
    wire [21:0] sum256_128_wire02  = {1'd0, sum512_256_wire03[20:0]}  + {1'd0, sum512_256_wire04[20:0]}  ;
    wire [21:0] sum256_128_wire03  = {1'd0, sum512_256_wire05[20:0]}  + {1'd0, sum512_256_wire06[20:0]}  ;
    wire [21:0] sum256_128_wire04  = {1'd0, sum512_256_wire07[20:0]}  + {1'd0, sum512_256_wire08[20:0]}  ;
    wire [21:0] sum256_128_wire05  = {1'd0, sum512_256_wire09[20:0]}  + {1'd0, sum512_256_wire10[20:0]}  ;
    wire [21:0] sum256_128_wire06  = {1'd0, sum512_256_wire11[20:0]}  + {1'd0, sum512_256_wire12[20:0]}  ;
    wire [21:0] sum256_128_wire07  = {1'd0, sum512_256_wire13[20:0]}  + {1'd0, sum512_256_wire14[20:0]}  ;
    wire [21:0] sum256_128_wire08  = {1'd0, sum512_256_wire15[20:0]}  + {1'd0, sum512_256_wire16[20:0]}  ;
    wire [21:0] sum256_128_wire09  = {1'd0, sum512_256_wire17[20:0]}  + {1'd0, sum512_256_wire18[20:0]}  ;
    wire [21:0] sum256_128_wire10  = {1'd0, sum512_256_wire19[20:0]}  + {1'd0, sum512_256_wire20[20:0]}  ;
    wire [21:0] sum256_128_wire11  = {1'd0, sum512_256_wire21[20:0]}  + {1'd0, sum512_256_wire22[20:0]}  ;
    wire [21:0] sum256_128_wire12  = {1'd0, sum512_256_wire23[20:0]}  + {1'd0, sum512_256_wire24[20:0]}  ;
    wire [21:0] sum256_128_wire13  = {1'd0, sum512_256_wire25[20:0]}  + {1'd0, sum512_256_wire26[20:0]}  ;
    wire [21:0] sum256_128_wire14  = {1'd0, sum512_256_wire27[20:0]}  + {1'd0, sum512_256_wire28[20:0]}  ;
    wire [21:0] sum256_128_wire15  = {1'd0, sum512_256_wire29[20:0]}  + {1'd0, sum512_256_wire30[20:0]}  ;
    wire [21:0] sum256_128_wire16  = {1'd0, sum512_256_wire31[20:0]}  + {1'd0, sum512_256_wire32[20:0]}  ;
    wire [21:0] sum256_128_wire17  = {1'd0, sum512_256_wire33[20:0]}  + {1'd0, sum512_256_wire34[20:0]}  ;
    wire [21:0] sum256_128_wire18  = {1'd0, sum512_256_wire35[20:0]}  + {1'd0, sum512_256_wire36[20:0]}  ;
    wire [21:0] sum256_128_wire19  = {1'd0, sum512_256_wire37[20:0]}  + {1'd0, sum512_256_wire38[20:0]}  ;
    wire [21:0] sum256_128_wire20  = {1'd0, sum512_256_wire39[20:0]}  + {1'd0, sum512_256_wire40[20:0]}  ;
    wire [21:0] sum256_128_wire21  = {1'd0, sum512_256_wire41[20:0]}  + {1'd0, sum512_256_wire42[20:0]}  ;
    wire [21:0] sum256_128_wire22  = {1'd0, sum512_256_wire43[20:0]}  + {1'd0, sum512_256_wire44[20:0]}  ;
    wire [21:0] sum256_128_wire23  = {1'd0, sum512_256_wire45[20:0]}  + {1'd0, sum512_256_wire46[20:0]}  ;
    wire [21:0] sum256_128_wire24  = {1'd0, sum512_256_wire47[20:0]}  + {1'd0, sum512_256_wire48[20:0]}  ;
    wire [21:0] sum256_128_wire25  = {1'd0, sum512_256_wire49[20:0]}  + {1'd0, sum512_256_wire50[20:0]}  ;
    wire [21:0] sum256_128_wire26  = {1'd0, sum512_256_wire51[20:0]}  + {1'd0, sum512_256_wire52[20:0]}  ;
    wire [21:0] sum256_128_wire27  = {1'd0, sum512_256_wire53[20:0]}  + {1'd0, sum512_256_wire54[20:0]}  ;
    wire [21:0] sum256_128_wire28  = {1'd0, sum512_256_wire55[20:0]}  + {1'd0, sum512_256_wire56[20:0]}  ;
    wire [21:0] sum256_128_wire29  = {1'd0, sum512_256_wire57[20:0]}  + {1'd0, sum512_256_wire58[20:0]}  ;
    wire [21:0] sum256_128_wire30  = {1'd0, sum512_256_wire59[20:0]}  + {1'd0, sum512_256_wire60[20:0]}  ;
    wire [21:0] sum256_128_wire31  = {1'd0, sum512_256_wire61[20:0]}  + {1'd0, sum512_256_wire62[20:0]}  ;
    wire [21:0] sum256_128_wire32  = {1'd0, sum512_256_wire63[20:0]}  + {1'd0, sum512_256_wire64[20:0]}  ;
    wire [21:0] sum256_128_wire33  = {1'd0, sum512_256_wire65[20:0]}  + {1'd0, sum512_256_wire66[20:0]}  ;
    wire [21:0] sum256_128_wire34  = {1'd0, sum512_256_wire67[20:0]}  + {1'd0, sum512_256_wire68[20:0]}  ;
    wire [21:0] sum256_128_wire35  = {1'd0, sum512_256_wire69[20:0]}  + {1'd0, sum512_256_wire70[20:0]}  ;
    wire [21:0] sum256_128_wire36  = {1'd0, sum512_256_wire71[20:0]}  + {1'd0, sum512_256_wire72[20:0]}  ;
    wire [21:0] sum256_128_wire37  = {1'd0, sum512_256_wire73[20:0]}  + {1'd0, sum512_256_wire74[20:0]}  ;
    wire [21:0] sum256_128_wire38  = {1'd0, sum512_256_wire75[20:0]}  + {1'd0, sum512_256_wire76[20:0]}  ;
    wire [21:0] sum256_128_wire39  = {1'd0, sum512_256_wire77[20:0]}  + {1'd0, sum512_256_wire78[20:0]}  ;
    wire [21:0] sum256_128_wire40  = {1'd0, sum512_256_wire79[20:0]}  + {1'd0, sum512_256_wire80[20:0]}  ;
    wire [21:0] sum256_128_wire41  = {1'd0, sum512_256_wire81[20:0]}  + {1'd0, sum512_256_wire82[20:0]}  ;
    wire [21:0] sum256_128_wire42  = {1'd0, sum512_256_wire83[20:0]}  + {1'd0, sum512_256_wire84[20:0]}  ;
    wire [21:0] sum256_128_wire43  = {1'd0, sum512_256_wire85[20:0]}  + {1'd0, sum512_256_wire86[20:0]}  ;
    wire [21:0] sum256_128_wire44  = {1'd0, sum512_256_wire87[20:0]}  + {1'd0, sum512_256_wire88[20:0]}  ;
    wire [21:0] sum256_128_wire45  = {1'd0, sum512_256_wire89[20:0]}  + {1'd0, sum512_256_wire90[20:0]}  ;
    wire [21:0] sum256_128_wire46  = {1'd0, sum512_256_wire91[20:0]}  + {1'd0, sum512_256_wire92[20:0]}  ;
    wire [21:0] sum256_128_wire47  = {1'd0, sum512_256_wire93[20:0]}  + {1'd0, sum512_256_wire94[20:0]}  ;
    wire [21:0] sum256_128_wire48  = {1'd0, sum512_256_wire95[20:0]}  + {1'd0, sum512_256_wire96[20:0]}  ;
    wire [21:0] sum256_128_wire49  = {1'd0, sum512_256_wire97[20:0]}  + {1'd0, sum512_256_wire98[20:0]}  ;
    wire [21:0] sum256_128_wire50  = {1'd0, sum512_256_wire99[20:0]}  + {1'd0, sum512_256_wire100[20:0]} ;
    wire [21:0] sum256_128_wire51  = {1'd0, sum512_256_wire101[20:0]} + {1'd0, sum512_256_wire102[20:0]} ;
    wire [21:0] sum256_128_wire52  = {1'd0, sum512_256_wire103[20:0]} + {1'd0, sum512_256_wire104[20:0]} ;
    wire [21:0] sum256_128_wire53  = {1'd0, sum512_256_wire105[20:0]} + {1'd0, sum512_256_wire106[20:0]} ;
    wire [21:0] sum256_128_wire54  = {1'd0, sum512_256_wire107[20:0]} + {1'd0, sum512_256_wire108[20:0]} ;
    wire [21:0] sum256_128_wire55  = {1'd0, sum512_256_wire109[20:0]} + {1'd0, sum512_256_wire110[20:0]} ;
    wire [21:0] sum256_128_wire56  = {1'd0, sum512_256_wire111[20:0]} + {1'd0, sum512_256_wire112[20:0]} ;
    wire [21:0] sum256_128_wire57  = {1'd0, sum512_256_wire113[20:0]} + {1'd0, sum512_256_wire114[20:0]} ;
    wire [21:0] sum256_128_wire58  = {1'd0, sum512_256_wire115[20:0]} + {1'd0, sum512_256_wire116[20:0]} ;
    wire [21:0] sum256_128_wire59  = {1'd0, sum512_256_wire117[20:0]} + {1'd0, sum512_256_wire118[20:0]} ;
    wire [21:0] sum256_128_wire60  = {1'd0, sum512_256_wire119[20:0]} + {1'd0, sum512_256_wire120[20:0]} ;
    wire [21:0] sum256_128_wire61  = {1'd0, sum512_256_wire121[20:0]} + {1'd0, sum512_256_wire122[20:0]} ;
    wire [21:0] sum256_128_wire62  = {1'd0, sum512_256_wire123[20:0]} + {1'd0, sum512_256_wire124[20:0]} ;
    wire [21:0] sum256_128_wire63  = {1'd0, sum512_256_wire125[20:0]} + {1'd0, sum512_256_wire126[20:0]} ;
    wire [21:0] sum256_128_wire64  = {1'd0, sum512_256_wire127[20:0]} + {1'd0, sum512_256_wire128[20:0]} ;
    wire [21:0] sum256_128_wire65  = {1'd0, sum512_256_wire129[20:0]} + {1'd0, sum512_256_wire130[20:0]} ;
    wire [21:0] sum256_128_wire66  = {1'd0, sum512_256_wire131[20:0]} + {1'd0, sum512_256_wire132[20:0]} ;
    wire [21:0] sum256_128_wire67  = {1'd0, sum512_256_wire133[20:0]} + {1'd0, sum512_256_wire134[20:0]} ;
    wire [21:0] sum256_128_wire68  = {1'd0, sum512_256_wire135[20:0]} + {1'd0, sum512_256_wire136[20:0]} ;
    wire [21:0] sum256_128_wire69  = {1'd0, sum512_256_wire137[20:0]} + {1'd0, sum512_256_wire138[20:0]} ;
    wire [21:0] sum256_128_wire70  = {1'd0, sum512_256_wire139[20:0]} + {1'd0, sum512_256_wire140[20:0]} ;
    wire [21:0] sum256_128_wire71  = {1'd0, sum512_256_wire141[20:0]} + {1'd0, sum512_256_wire142[20:0]} ;
    wire [21:0] sum256_128_wire72  = {1'd0, sum512_256_wire143[20:0]} + {1'd0, sum512_256_wire144[20:0]} ;
    wire [21:0] sum256_128_wire73  = {1'd0, sum512_256_wire145[20:0]} + {1'd0, sum512_256_wire146[20:0]} ;
    wire [21:0] sum256_128_wire74  = {1'd0, sum512_256_wire147[20:0]} + {1'd0, sum512_256_wire148[20:0]} ;
    wire [21:0] sum256_128_wire75  = {1'd0, sum512_256_wire149[20:0]} + {1'd0, sum512_256_wire150[20:0]} ;
    wire [21:0] sum256_128_wire76  = {1'd0, sum512_256_wire151[20:0]} + {1'd0, sum512_256_wire152[20:0]} ;
    wire [21:0] sum256_128_wire77  = {1'd0, sum512_256_wire153[20:0]} + {1'd0, sum512_256_wire154[20:0]} ;
    wire [21:0] sum256_128_wire78  = {1'd0, sum512_256_wire155[20:0]} + {1'd0, sum512_256_wire156[20:0]} ;
    wire [21:0] sum256_128_wire79  = {1'd0, sum512_256_wire157[20:0]} + {1'd0, sum512_256_wire158[20:0]} ;
    wire [21:0] sum256_128_wire80  = {1'd0, sum512_256_wire159[20:0]} + {1'd0, sum512_256_wire160[20:0]} ;
    wire [21:0] sum256_128_wire81  = {1'd0, sum512_256_wire161[20:0]} + {1'd0, sum512_256_wire162[20:0]} ;
    wire [21:0] sum256_128_wire82  = {1'd0, sum512_256_wire163[20:0]} + {1'd0, sum512_256_wire164[20:0]} ;
    wire [21:0] sum256_128_wire83  = {1'd0, sum512_256_wire165[20:0]} + {1'd0, sum512_256_wire166[20:0]} ;
    wire [21:0] sum256_128_wire84  = {1'd0, sum512_256_wire167[20:0]} + {1'd0, sum512_256_wire168[20:0]} ;
    wire [21:0] sum256_128_wire85  = {1'd0, sum512_256_wire169[20:0]} + {1'd0, sum512_256_wire170[20:0]} ;
    wire [21:0] sum256_128_wire86  = {1'd0, sum512_256_wire171[20:0]} + {1'd0, sum512_256_wire172[20:0]} ;
    wire [21:0] sum256_128_wire87  = {1'd0, sum512_256_wire173[20:0]} + {1'd0, sum512_256_wire174[20:0]} ;
    wire [21:0] sum256_128_wire88  = {1'd0, sum512_256_wire175[20:0]} + {1'd0, sum512_256_wire176[20:0]} ;
    wire [21:0] sum256_128_wire89  = {1'd0, sum512_256_wire177[20:0]} + {1'd0, sum512_256_wire178[20:0]} ;
    wire [21:0] sum256_128_wire90  = {1'd0, sum512_256_wire179[20:0]} + {1'd0, sum512_256_wire180[20:0]} ;
    wire [21:0] sum256_128_wire91  = {1'd0, sum512_256_wire181[20:0]} + {1'd0, sum512_256_wire182[20:0]} ;
    wire [21:0] sum256_128_wire92  = {1'd0, sum512_256_wire183[20:0]} + {1'd0, sum512_256_wire184[20:0]} ;
    wire [21:0] sum256_128_wire93  = {1'd0, sum512_256_wire185[20:0]} + {1'd0, sum512_256_wire186[20:0]} ;
    wire [21:0] sum256_128_wire94  = {1'd0, sum512_256_wire187[20:0]} + {1'd0, sum512_256_wire188[20:0]} ;
    wire [21:0] sum256_128_wire95  = {1'd0, sum512_256_wire189[20:0]} + {1'd0, sum512_256_wire190[20:0]} ;
    wire [21:0] sum256_128_wire96  = {1'd0, sum512_256_wire191[20:0]} + {1'd0, sum512_256_wire192[20:0]} ;
    wire [21:0] sum256_128_wire97  = {1'd0, sum512_256_wire193[20:0]} + {1'd0, sum512_256_wire194[20:0]} ;
    wire [21:0] sum256_128_wire98  = {1'd0, sum512_256_wire195[20:0]} + {1'd0, sum512_256_wire196[20:0]} ;
    wire [21:0] sum256_128_wire99  = {1'd0, sum512_256_wire197[20:0]} + {1'd0, sum512_256_wire198[20:0]} ;
    wire [21:0] sum256_128_wire100 = {1'd0, sum512_256_wire199[20:0]} + {1'd0, sum512_256_wire200[20:0]} ;
    wire [21:0] sum256_128_wire101 = {1'd0, sum512_256_wire201[20:0]} + {1'd0, sum512_256_wire202[20:0]} ;
    wire [21:0] sum256_128_wire102 = {1'd0, sum512_256_wire203[20:0]} + {1'd0, sum512_256_wire204[20:0]} ;
    wire [21:0] sum256_128_wire103 = {1'd0, sum512_256_wire205[20:0]} + {1'd0, sum512_256_wire206[20:0]} ;
    wire [21:0] sum256_128_wire104 = {1'd0, sum512_256_wire207[20:0]} + {1'd0, sum512_256_wire208[20:0]} ;
    wire [21:0] sum256_128_wire105 = {1'd0, sum512_256_wire209[20:0]} + {1'd0, sum512_256_wire210[20:0]} ;
    wire [21:0] sum256_128_wire106 = {1'd0, sum512_256_wire211[20:0]} + {1'd0, sum512_256_wire212[20:0]} ;
    wire [21:0] sum256_128_wire107 = {1'd0, sum512_256_wire213[20:0]} + {1'd0, sum512_256_wire214[20:0]} ;
    wire [21:0] sum256_128_wire108 = {1'd0, sum512_256_wire215[20:0]} + {1'd0, sum512_256_wire216[20:0]} ;
    wire [21:0] sum256_128_wire109 = {1'd0, sum512_256_wire217[20:0]} + {1'd0, sum512_256_wire218[20:0]} ;
    wire [21:0] sum256_128_wire110 = {1'd0, sum512_256_wire219[20:0]} + {1'd0, sum512_256_wire220[20:0]} ;
    wire [21:0] sum256_128_wire111 = {1'd0, sum512_256_wire221[20:0]} + {1'd0, sum512_256_wire222[20:0]} ;
    wire [21:0] sum256_128_wire112 = {1'd0, sum512_256_wire223[20:0]} + {1'd0, sum512_256_wire224[20:0]} ;
    wire [21:0] sum256_128_wire113 = {1'd0, sum512_256_wire225[20:0]} + {1'd0, sum512_256_wire226[20:0]} ;
    wire [21:0] sum256_128_wire114 = {1'd0, sum512_256_wire227[20:0]} + {1'd0, sum512_256_wire228[20:0]} ;
    wire [21:0] sum256_128_wire115 = {1'd0, sum512_256_wire229[20:0]} + {1'd0, sum512_256_wire230[20:0]} ;
    wire [21:0] sum256_128_wire116 = {1'd0, sum512_256_wire231[20:0]} + {1'd0, sum512_256_wire232[20:0]} ;
    wire [21:0] sum256_128_wire117 = {1'd0, sum512_256_wire233[20:0]} + {1'd0, sum512_256_wire234[20:0]} ;
    wire [21:0] sum256_128_wire118 = {1'd0, sum512_256_wire235[20:0]} + {1'd0, sum512_256_wire236[20:0]} ;
    wire [21:0] sum256_128_wire119 = {1'd0, sum512_256_wire237[20:0]} + {1'd0, sum512_256_wire238[20:0]} ;
    wire [21:0] sum256_128_wire120 = {1'd0, sum512_256_wire239[20:0]} + {1'd0, sum512_256_wire240[20:0]} ;
    wire [21:0] sum256_128_wire121 = {1'd0, sum512_256_wire241[20:0]} + {1'd0, sum512_256_wire242[20:0]} ;
    wire [21:0] sum256_128_wire122 = {1'd0, sum512_256_wire243[20:0]} + {1'd0, sum512_256_wire244[20:0]} ;
    wire [21:0] sum256_128_wire123 = {1'd0, sum512_256_wire245[20:0]} + {1'd0, sum512_256_wire246[20:0]} ;
    wire [21:0] sum256_128_wire124 = {1'd0, sum512_256_wire247[20:0]} + {1'd0, sum512_256_wire248[20:0]} ;
    wire [21:0] sum256_128_wire125 = {1'd0, sum512_256_wire249[20:0]} + {1'd0, sum512_256_wire250[20:0]} ;
    wire [21:0] sum256_128_wire126 = {1'd0, sum512_256_wire251[20:0]} + {1'd0, sum512_256_wire252[20:0]} ;
    wire [21:0] sum256_128_wire127 = {1'd0, sum512_256_wire253[20:0]} + {1'd0, sum512_256_wire254[20:0]} ;
    wire [21:0] sum256_128_wire128 = {1'd0, sum512_256_wire255[20:0]} + {1'd0, sum512_256_wire256[20:0]} ;
   
    reg [21:0] sum256_128_reg01,  sum256_128_reg02,  sum256_128_reg03,  sum256_128_reg04,
               sum256_128_reg05,  sum256_128_reg06,  sum256_128_reg07,  sum256_128_reg08,
               sum256_128_reg09,  sum256_128_reg10,  sum256_128_reg11,  sum256_128_reg12,
               sum256_128_reg13,  sum256_128_reg14,  sum256_128_reg15,  sum256_128_reg16,
               sum256_128_reg17,  sum256_128_reg18,  sum256_128_reg19,  sum256_128_reg20,
               sum256_128_reg21,  sum256_128_reg22,  sum256_128_reg23,  sum256_128_reg24,
               sum256_128_reg25,  sum256_128_reg26,  sum256_128_reg27,  sum256_128_reg28,
               sum256_128_reg29,  sum256_128_reg30,  sum256_128_reg31,  sum256_128_reg32,
               sum256_128_reg33,  sum256_128_reg34,  sum256_128_reg35,  sum256_128_reg36,
               sum256_128_reg37,  sum256_128_reg38,  sum256_128_reg39,  sum256_128_reg40,
               sum256_128_reg41,  sum256_128_reg42,  sum256_128_reg43,  sum256_128_reg44,
               sum256_128_reg45,  sum256_128_reg46,  sum256_128_reg47,  sum256_128_reg48,
               sum256_128_reg49,  sum256_128_reg50,  sum256_128_reg51,  sum256_128_reg52,
               sum256_128_reg53,  sum256_128_reg54,  sum256_128_reg55,  sum256_128_reg56,
               sum256_128_reg57,  sum256_128_reg58,  sum256_128_reg59,  sum256_128_reg60,
               sum256_128_reg61,  sum256_128_reg62,  sum256_128_reg63,  sum256_128_reg64,
               sum256_128_reg65,  sum256_128_reg66,  sum256_128_reg67,  sum256_128_reg68,
               sum256_128_reg69,  sum256_128_reg70,  sum256_128_reg71,  sum256_128_reg72,
               sum256_128_reg73,  sum256_128_reg74,  sum256_128_reg75,  sum256_128_reg76,
               sum256_128_reg77,  sum256_128_reg78,  sum256_128_reg79,  sum256_128_reg80,
               sum256_128_reg81,  sum256_128_reg82,  sum256_128_reg83,  sum256_128_reg84,
               sum256_128_reg85,  sum256_128_reg86,  sum256_128_reg87,  sum256_128_reg88,
               sum256_128_reg89,  sum256_128_reg90,  sum256_128_reg91,  sum256_128_reg92,
               sum256_128_reg93,  sum256_128_reg94,  sum256_128_reg95,  sum256_128_reg96,
               sum256_128_reg97,  sum256_128_reg98,  sum256_128_reg99,  sum256_128_reg100,
               sum256_128_reg101, sum256_128_reg102, sum256_128_reg103, sum256_128_reg104,
               sum256_128_reg105, sum256_128_reg106, sum256_128_reg107, sum256_128_reg108,
               sum256_128_reg109, sum256_128_reg110, sum256_128_reg111, sum256_128_reg112,
               sum256_128_reg113, sum256_128_reg114, sum256_128_reg115, sum256_128_reg116,
               sum256_128_reg117, sum256_128_reg118, sum256_128_reg119, sum256_128_reg120,
               sum256_128_reg121, sum256_128_reg122, sum256_128_reg123, sum256_128_reg124,
               sum256_128_reg125, sum256_128_reg126, sum256_128_reg127, sum256_128_reg128;

    always @ (posedge clk) begin
		if(rst) begin
            sum256_128_reg01[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg02[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg03[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg04[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg05[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg06[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg07[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg08[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg09[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg10[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg11[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg12[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg13[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg14[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg15[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg16[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg17[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg18[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg19[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg20[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg21[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg22[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg23[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg24[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg25[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg26[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg27[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg28[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg29[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg30[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg31[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg32[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg33[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg34[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg35[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg36[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg37[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg38[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg39[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg40[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg41[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg42[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg43[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg44[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg45[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg46[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg47[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg48[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg49[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg50[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg51[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg52[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg53[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg54[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg55[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg56[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg57[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg58[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg59[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg60[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg61[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg62[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg63[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg64[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg65[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg66[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg67[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg68[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg69[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg70[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg71[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg72[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg73[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg74[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg75[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg76[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg77[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg78[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg79[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg80[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg81[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg82[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg83[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg84[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg85[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg86[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg87[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg88[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg89[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg90[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg91[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg92[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg93[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg94[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg95[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg96[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg97[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg98[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg99[21:0]  <= #DLY 22'd0 ;
            sum256_128_reg100[21:0] <= #DLY 22'd0 ;
            sum256_128_reg101[21:0] <= #DLY 22'd0 ;
            sum256_128_reg102[21:0] <= #DLY 22'd0 ;
            sum256_128_reg103[21:0] <= #DLY 22'd0 ;
            sum256_128_reg104[21:0] <= #DLY 22'd0 ;
            sum256_128_reg105[21:0] <= #DLY 22'd0 ;
            sum256_128_reg106[21:0] <= #DLY 22'd0 ;
            sum256_128_reg107[21:0] <= #DLY 22'd0 ;
            sum256_128_reg108[21:0] <= #DLY 22'd0 ;
            sum256_128_reg109[21:0] <= #DLY 22'd0 ;
            sum256_128_reg110[21:0] <= #DLY 22'd0 ;
            sum256_128_reg111[21:0] <= #DLY 22'd0 ;
            sum256_128_reg112[21:0] <= #DLY 22'd0 ;
            sum256_128_reg113[21:0] <= #DLY 22'd0 ;
            sum256_128_reg114[21:0] <= #DLY 22'd0 ;
            sum256_128_reg115[21:0] <= #DLY 22'd0 ;
            sum256_128_reg116[21:0] <= #DLY 22'd0 ;
            sum256_128_reg117[21:0] <= #DLY 22'd0 ;
            sum256_128_reg118[21:0] <= #DLY 22'd0 ;
            sum256_128_reg119[21:0] <= #DLY 22'd0 ;
            sum256_128_reg120[21:0] <= #DLY 22'd0 ;
            sum256_128_reg121[21:0] <= #DLY 22'd0 ;
            sum256_128_reg122[21:0] <= #DLY 22'd0 ;
            sum256_128_reg123[21:0] <= #DLY 22'd0 ;
            sum256_128_reg124[21:0] <= #DLY 22'd0 ;
            sum256_128_reg125[21:0] <= #DLY 22'd0 ;
            sum256_128_reg126[21:0] <= #DLY 22'd0 ;
            sum256_128_reg127[21:0] <= #DLY 22'd0 ;
            sum256_128_reg128[21:0] <= #DLY 22'd0 ;
		end else begin
            sum256_128_reg01[21:0]  <= #DLY sum256_128_wire01[21:0]  ;
            sum256_128_reg02[21:0]  <= #DLY sum256_128_wire02[21:0]  ;
            sum256_128_reg03[21:0]  <= #DLY sum256_128_wire03[21:0]  ;
            sum256_128_reg04[21:0]  <= #DLY sum256_128_wire04[21:0]  ;
            sum256_128_reg05[21:0]  <= #DLY sum256_128_wire05[21:0]  ;
            sum256_128_reg06[21:0]  <= #DLY sum256_128_wire06[21:0]  ;
            sum256_128_reg07[21:0]  <= #DLY sum256_128_wire07[21:0]  ;
            sum256_128_reg08[21:0]  <= #DLY sum256_128_wire08[21:0]  ;
            sum256_128_reg09[21:0]  <= #DLY sum256_128_wire09[21:0]  ;
            sum256_128_reg10[21:0]  <= #DLY sum256_128_wire10[21:0]  ;
            sum256_128_reg11[21:0]  <= #DLY sum256_128_wire11[21:0]  ;
            sum256_128_reg12[21:0]  <= #DLY sum256_128_wire12[21:0]  ;
            sum256_128_reg13[21:0]  <= #DLY sum256_128_wire13[21:0]  ;
            sum256_128_reg14[21:0]  <= #DLY sum256_128_wire14[21:0]  ;
            sum256_128_reg15[21:0]  <= #DLY sum256_128_wire15[21:0]  ;
            sum256_128_reg16[21:0]  <= #DLY sum256_128_wire16[21:0]  ;
            sum256_128_reg17[21:0]  <= #DLY sum256_128_wire17[21:0]  ;
            sum256_128_reg18[21:0]  <= #DLY sum256_128_wire18[21:0]  ;
            sum256_128_reg19[21:0]  <= #DLY sum256_128_wire19[21:0]  ;
            sum256_128_reg20[21:0]  <= #DLY sum256_128_wire20[21:0]  ;
            sum256_128_reg21[21:0]  <= #DLY sum256_128_wire21[21:0]  ;
            sum256_128_reg22[21:0]  <= #DLY sum256_128_wire22[21:0]  ;
            sum256_128_reg23[21:0]  <= #DLY sum256_128_wire23[21:0]  ;
            sum256_128_reg24[21:0]  <= #DLY sum256_128_wire24[21:0]  ;
            sum256_128_reg25[21:0]  <= #DLY sum256_128_wire25[21:0]  ;
            sum256_128_reg26[21:0]  <= #DLY sum256_128_wire26[21:0]  ;
            sum256_128_reg27[21:0]  <= #DLY sum256_128_wire27[21:0]  ;
            sum256_128_reg28[21:0]  <= #DLY sum256_128_wire28[21:0]  ;
            sum256_128_reg29[21:0]  <= #DLY sum256_128_wire29[21:0]  ;
            sum256_128_reg30[21:0]  <= #DLY sum256_128_wire30[21:0]  ;
            sum256_128_reg31[21:0]  <= #DLY sum256_128_wire31[21:0]  ;
            sum256_128_reg32[21:0]  <= #DLY sum256_128_wire32[21:0]  ;
            sum256_128_reg33[21:0]  <= #DLY sum256_128_wire33[21:0]  ;
            sum256_128_reg34[21:0]  <= #DLY sum256_128_wire34[21:0]  ;
            sum256_128_reg35[21:0]  <= #DLY sum256_128_wire35[21:0]  ;
            sum256_128_reg36[21:0]  <= #DLY sum256_128_wire36[21:0]  ;
            sum256_128_reg37[21:0]  <= #DLY sum256_128_wire37[21:0]  ;
            sum256_128_reg38[21:0]  <= #DLY sum256_128_wire38[21:0]  ;
            sum256_128_reg39[21:0]  <= #DLY sum256_128_wire39[21:0]  ;
            sum256_128_reg40[21:0]  <= #DLY sum256_128_wire40[21:0]  ;
            sum256_128_reg41[21:0]  <= #DLY sum256_128_wire41[21:0]  ;
            sum256_128_reg42[21:0]  <= #DLY sum256_128_wire42[21:0]  ;
            sum256_128_reg43[21:0]  <= #DLY sum256_128_wire43[21:0]  ;
            sum256_128_reg44[21:0]  <= #DLY sum256_128_wire44[21:0]  ;
            sum256_128_reg45[21:0]  <= #DLY sum256_128_wire45[21:0]  ;
            sum256_128_reg46[21:0]  <= #DLY sum256_128_wire46[21:0]  ;
            sum256_128_reg47[21:0]  <= #DLY sum256_128_wire47[21:0]  ;
            sum256_128_reg48[21:0]  <= #DLY sum256_128_wire48[21:0]  ;
            sum256_128_reg49[21:0]  <= #DLY sum256_128_wire49[21:0]  ;
            sum256_128_reg50[21:0]  <= #DLY sum256_128_wire50[21:0]  ;
            sum256_128_reg51[21:0]  <= #DLY sum256_128_wire51[21:0]  ;
            sum256_128_reg52[21:0]  <= #DLY sum256_128_wire52[21:0]  ;
            sum256_128_reg53[21:0]  <= #DLY sum256_128_wire53[21:0]  ;
            sum256_128_reg54[21:0]  <= #DLY sum256_128_wire54[21:0]  ;
            sum256_128_reg55[21:0]  <= #DLY sum256_128_wire55[21:0]  ;
            sum256_128_reg56[21:0]  <= #DLY sum256_128_wire56[21:0]  ;
            sum256_128_reg57[21:0]  <= #DLY sum256_128_wire57[21:0]  ;
            sum256_128_reg58[21:0]  <= #DLY sum256_128_wire58[21:0]  ;
            sum256_128_reg59[21:0]  <= #DLY sum256_128_wire59[21:0]  ;
            sum256_128_reg60[21:0]  <= #DLY sum256_128_wire60[21:0]  ;
            sum256_128_reg61[21:0]  <= #DLY sum256_128_wire61[21:0]  ;
            sum256_128_reg62[21:0]  <= #DLY sum256_128_wire62[21:0]  ;
            sum256_128_reg63[21:0]  <= #DLY sum256_128_wire63[21:0]  ;
            sum256_128_reg64[21:0]  <= #DLY sum256_128_wire64[21:0]  ;
            sum256_128_reg65[21:0]  <= #DLY sum256_128_wire65[21:0]  ;
            sum256_128_reg66[21:0]  <= #DLY sum256_128_wire66[21:0]  ;
            sum256_128_reg67[21:0]  <= #DLY sum256_128_wire67[21:0]  ;
            sum256_128_reg68[21:0]  <= #DLY sum256_128_wire68[21:0]  ;
            sum256_128_reg69[21:0]  <= #DLY sum256_128_wire69[21:0]  ;
            sum256_128_reg70[21:0]  <= #DLY sum256_128_wire70[21:0]  ;
            sum256_128_reg71[21:0]  <= #DLY sum256_128_wire71[21:0]  ;
            sum256_128_reg72[21:0]  <= #DLY sum256_128_wire72[21:0]  ;
            sum256_128_reg73[21:0]  <= #DLY sum256_128_wire73[21:0]  ;
            sum256_128_reg74[21:0]  <= #DLY sum256_128_wire74[21:0]  ;
            sum256_128_reg75[21:0]  <= #DLY sum256_128_wire75[21:0]  ;
            sum256_128_reg76[21:0]  <= #DLY sum256_128_wire76[21:0]  ;
            sum256_128_reg77[21:0]  <= #DLY sum256_128_wire77[21:0]  ;
            sum256_128_reg78[21:0]  <= #DLY sum256_128_wire78[21:0]  ;
            sum256_128_reg79[21:0]  <= #DLY sum256_128_wire79[21:0]  ;
            sum256_128_reg80[21:0]  <= #DLY sum256_128_wire80[21:0]  ;
            sum256_128_reg81[21:0]  <= #DLY sum256_128_wire81[21:0]  ;
            sum256_128_reg82[21:0]  <= #DLY sum256_128_wire82[21:0]  ;
            sum256_128_reg83[21:0]  <= #DLY sum256_128_wire83[21:0]  ;
            sum256_128_reg84[21:0]  <= #DLY sum256_128_wire84[21:0]  ;
            sum256_128_reg85[21:0]  <= #DLY sum256_128_wire85[21:0]  ;
            sum256_128_reg86[21:0]  <= #DLY sum256_128_wire86[21:0]  ;
            sum256_128_reg87[21:0]  <= #DLY sum256_128_wire87[21:0]  ;
            sum256_128_reg88[21:0]  <= #DLY sum256_128_wire88[21:0]  ;
            sum256_128_reg89[21:0]  <= #DLY sum256_128_wire89[21:0]  ;
            sum256_128_reg90[21:0]  <= #DLY sum256_128_wire90[21:0]  ;
            sum256_128_reg91[21:0]  <= #DLY sum256_128_wire91[21:0]  ;
            sum256_128_reg92[21:0]  <= #DLY sum256_128_wire92[21:0]  ;
            sum256_128_reg93[21:0]  <= #DLY sum256_128_wire93[21:0]  ;
            sum256_128_reg94[21:0]  <= #DLY sum256_128_wire94[21:0]  ;
            sum256_128_reg95[21:0]  <= #DLY sum256_128_wire95[21:0]  ;
            sum256_128_reg96[21:0]  <= #DLY sum256_128_wire96[21:0]  ;
            sum256_128_reg97[21:0]  <= #DLY sum256_128_wire97[21:0]  ;
            sum256_128_reg98[21:0]  <= #DLY sum256_128_wire98[21:0]  ;
            sum256_128_reg99[21:0]  <= #DLY sum256_128_wire99[21:0]  ;
            sum256_128_reg100[21:0] <= #DLY sum256_128_wire100[21:0] ;
            sum256_128_reg101[21:0] <= #DLY sum256_128_wire101[21:0] ;
            sum256_128_reg102[21:0] <= #DLY sum256_128_wire102[21:0] ;
            sum256_128_reg103[21:0] <= #DLY sum256_128_wire103[21:0] ;
            sum256_128_reg104[21:0] <= #DLY sum256_128_wire104[21:0] ;
            sum256_128_reg105[21:0] <= #DLY sum256_128_wire105[21:0] ;
            sum256_128_reg106[21:0] <= #DLY sum256_128_wire106[21:0] ;
            sum256_128_reg107[21:0] <= #DLY sum256_128_wire107[21:0] ;
            sum256_128_reg108[21:0] <= #DLY sum256_128_wire108[21:0] ;
            sum256_128_reg109[21:0] <= #DLY sum256_128_wire109[21:0] ;
            sum256_128_reg110[21:0] <= #DLY sum256_128_wire110[21:0] ;
            sum256_128_reg111[21:0] <= #DLY sum256_128_wire111[21:0] ;
            sum256_128_reg112[21:0] <= #DLY sum256_128_wire112[21:0] ;
            sum256_128_reg113[21:0] <= #DLY sum256_128_wire113[21:0] ;
            sum256_128_reg114[21:0] <= #DLY sum256_128_wire114[21:0] ;
            sum256_128_reg115[21:0] <= #DLY sum256_128_wire115[21:0] ;
            sum256_128_reg116[21:0] <= #DLY sum256_128_wire116[21:0] ;
            sum256_128_reg117[21:0] <= #DLY sum256_128_wire117[21:0] ;
            sum256_128_reg118[21:0] <= #DLY sum256_128_wire118[21:0] ;
            sum256_128_reg119[21:0] <= #DLY sum256_128_wire119[21:0] ;
            sum256_128_reg120[21:0] <= #DLY sum256_128_wire120[21:0] ;
            sum256_128_reg121[21:0] <= #DLY sum256_128_wire121[21:0] ;
            sum256_128_reg122[21:0] <= #DLY sum256_128_wire122[21:0] ;
            sum256_128_reg123[21:0] <= #DLY sum256_128_wire123[21:0] ;
            sum256_128_reg124[21:0] <= #DLY sum256_128_wire124[21:0] ;
            sum256_128_reg125[21:0] <= #DLY sum256_128_wire125[21:0] ;
            sum256_128_reg126[21:0] <= #DLY sum256_128_wire126[21:0] ;
            sum256_128_reg127[21:0] <= #DLY sum256_128_wire127[21:0] ;
            sum256_128_reg128[21:0] <= #DLY sum256_128_wire128[21:0] ;
		end
	end
//
    /****************************
    // pipeline[35] Active
    ****************************/
    wire [22:0] sum128_64_wire01  = {1'd0, sum256_128_reg01[21:0]}  + {1'd0, sum256_128_reg02[21:0]}  ;
    wire [22:0] sum128_64_wire02  = {1'd0, sum256_128_reg03[21:0]}  + {1'd0, sum256_128_reg04[21:0]}  ;
    wire [22:0] sum128_64_wire03  = {1'd0, sum256_128_reg05[21:0]}  + {1'd0, sum256_128_reg06[21:0]}  ;
    wire [22:0] sum128_64_wire04  = {1'd0, sum256_128_reg07[21:0]}  + {1'd0, sum256_128_reg08[21:0]}  ;
    wire [22:0] sum128_64_wire05  = {1'd0, sum256_128_reg09[21:0]}  + {1'd0, sum256_128_reg10[21:0]}  ;
    wire [22:0] sum128_64_wire06  = {1'd0, sum256_128_reg11[21:0]}  + {1'd0, sum256_128_reg12[21:0]}  ;
    wire [22:0] sum128_64_wire07  = {1'd0, sum256_128_reg13[21:0]}  + {1'd0, sum256_128_reg14[21:0]}  ;
    wire [22:0] sum128_64_wire08  = {1'd0, sum256_128_reg15[21:0]}  + {1'd0, sum256_128_reg16[21:0]}  ;
    wire [22:0] sum128_64_wire09  = {1'd0, sum256_128_reg17[21:0]}  + {1'd0, sum256_128_reg18[21:0]}  ;
    wire [22:0] sum128_64_wire10  = {1'd0, sum256_128_reg19[21:0]}  + {1'd0, sum256_128_reg20[21:0]}  ;
    wire [22:0] sum128_64_wire11  = {1'd0, sum256_128_reg21[21:0]}  + {1'd0, sum256_128_reg22[21:0]}  ;
    wire [22:0] sum128_64_wire12  = {1'd0, sum256_128_reg23[21:0]}  + {1'd0, sum256_128_reg24[21:0]}  ;
    wire [22:0] sum128_64_wire13  = {1'd0, sum256_128_reg25[21:0]}  + {1'd0, sum256_128_reg26[21:0]}  ;
    wire [22:0] sum128_64_wire14  = {1'd0, sum256_128_reg27[21:0]}  + {1'd0, sum256_128_reg28[21:0]}  ;
    wire [22:0] sum128_64_wire15  = {1'd0, sum256_128_reg29[21:0]}  + {1'd0, sum256_128_reg30[21:0]}  ;
    wire [22:0] sum128_64_wire16  = {1'd0, sum256_128_reg31[21:0]}  + {1'd0, sum256_128_reg32[21:0]}  ;
    wire [22:0] sum128_64_wire17  = {1'd0, sum256_128_reg33[21:0]}  + {1'd0, sum256_128_reg34[21:0]}  ;
    wire [22:0] sum128_64_wire18  = {1'd0, sum256_128_reg35[21:0]}  + {1'd0, sum256_128_reg36[21:0]}  ;
    wire [22:0] sum128_64_wire19  = {1'd0, sum256_128_reg37[21:0]}  + {1'd0, sum256_128_reg38[21:0]}  ;
    wire [22:0] sum128_64_wire20  = {1'd0, sum256_128_reg39[21:0]}  + {1'd0, sum256_128_reg40[21:0]}  ;
    wire [22:0] sum128_64_wire21  = {1'd0, sum256_128_reg41[21:0]}  + {1'd0, sum256_128_reg42[21:0]}  ;
    wire [22:0] sum128_64_wire22  = {1'd0, sum256_128_reg43[21:0]}  + {1'd0, sum256_128_reg44[21:0]}  ;
    wire [22:0] sum128_64_wire23  = {1'd0, sum256_128_reg45[21:0]}  + {1'd0, sum256_128_reg46[21:0]}  ;
    wire [22:0] sum128_64_wire24  = {1'd0, sum256_128_reg47[21:0]}  + {1'd0, sum256_128_reg48[21:0]}  ;
    wire [22:0] sum128_64_wire25  = {1'd0, sum256_128_reg49[21:0]}  + {1'd0, sum256_128_reg50[21:0]}  ;
    wire [22:0] sum128_64_wire26  = {1'd0, sum256_128_reg51[21:0]}  + {1'd0, sum256_128_reg52[21:0]}  ;
    wire [22:0] sum128_64_wire27  = {1'd0, sum256_128_reg53[21:0]}  + {1'd0, sum256_128_reg54[21:0]}  ;
    wire [22:0] sum128_64_wire28  = {1'd0, sum256_128_reg55[21:0]}  + {1'd0, sum256_128_reg56[21:0]}  ;
    wire [22:0] sum128_64_wire29  = {1'd0, sum256_128_reg57[21:0]}  + {1'd0, sum256_128_reg58[21:0]}  ;
    wire [22:0] sum128_64_wire30  = {1'd0, sum256_128_reg59[21:0]}  + {1'd0, sum256_128_reg60[21:0]}  ;
    wire [22:0] sum128_64_wire31  = {1'd0, sum256_128_reg61[21:0]}  + {1'd0, sum256_128_reg62[21:0]}  ;
    wire [22:0] sum128_64_wire32  = {1'd0, sum256_128_reg63[21:0]}  + {1'd0, sum256_128_reg64[21:0]}  ;
    wire [22:0] sum128_64_wire33  = {1'd0, sum256_128_reg65[21:0]}  + {1'd0, sum256_128_reg66[21:0]}  ;
    wire [22:0] sum128_64_wire34  = {1'd0, sum256_128_reg67[21:0]}  + {1'd0, sum256_128_reg68[21:0]}  ;
    wire [22:0] sum128_64_wire35  = {1'd0, sum256_128_reg69[21:0]}  + {1'd0, sum256_128_reg70[21:0]}  ;
    wire [22:0] sum128_64_wire36  = {1'd0, sum256_128_reg71[21:0]}  + {1'd0, sum256_128_reg72[21:0]}  ;
    wire [22:0] sum128_64_wire37  = {1'd0, sum256_128_reg73[21:0]}  + {1'd0, sum256_128_reg74[21:0]}  ;
    wire [22:0] sum128_64_wire38  = {1'd0, sum256_128_reg75[21:0]}  + {1'd0, sum256_128_reg76[21:0]}  ;
    wire [22:0] sum128_64_wire39  = {1'd0, sum256_128_reg77[21:0]}  + {1'd0, sum256_128_reg78[21:0]}  ;
    wire [22:0] sum128_64_wire40  = {1'd0, sum256_128_reg79[21:0]}  + {1'd0, sum256_128_reg80[21:0]}  ;
    wire [22:0] sum128_64_wire41  = {1'd0, sum256_128_reg81[21:0]}  + {1'd0, sum256_128_reg82[21:0]}  ;
    wire [22:0] sum128_64_wire42  = {1'd0, sum256_128_reg83[21:0]}  + {1'd0, sum256_128_reg84[21:0]}  ;
    wire [22:0] sum128_64_wire43  = {1'd0, sum256_128_reg85[21:0]}  + {1'd0, sum256_128_reg86[21:0]}  ;
    wire [22:0] sum128_64_wire44  = {1'd0, sum256_128_reg87[21:0]}  + {1'd0, sum256_128_reg88[21:0]}  ;
    wire [22:0] sum128_64_wire45  = {1'd0, sum256_128_reg89[21:0]}  + {1'd0, sum256_128_reg90[21:0]}  ;
    wire [22:0] sum128_64_wire46  = {1'd0, sum256_128_reg91[21:0]}  + {1'd0, sum256_128_reg92[21:0]}  ;
    wire [22:0] sum128_64_wire47  = {1'd0, sum256_128_reg93[21:0]}  + {1'd0, sum256_128_reg94[21:0]}  ;
    wire [22:0] sum128_64_wire48  = {1'd0, sum256_128_reg95[21:0]}  + {1'd0, sum256_128_reg96[21:0]}  ;
    wire [22:0] sum128_64_wire49  = {1'd0, sum256_128_reg97[21:0]}  + {1'd0, sum256_128_reg98[21:0]}  ;
    wire [22:0] sum128_64_wire50  = {1'd0, sum256_128_reg99[21:0]}  + {1'd0, sum256_128_reg100[21:0]} ;
    wire [22:0] sum128_64_wire51  = {1'd0, sum256_128_reg101[21:0]} + {1'd0, sum256_128_reg102[21:0]} ;
    wire [22:0] sum128_64_wire52  = {1'd0, sum256_128_reg103[21:0]} + {1'd0, sum256_128_reg104[21:0]} ;
    wire [22:0] sum128_64_wire53  = {1'd0, sum256_128_reg105[21:0]} + {1'd0, sum256_128_reg106[21:0]} ;
    wire [22:0] sum128_64_wire54  = {1'd0, sum256_128_reg107[21:0]} + {1'd0, sum256_128_reg108[21:0]} ;
    wire [22:0] sum128_64_wire55  = {1'd0, sum256_128_reg109[21:0]} + {1'd0, sum256_128_reg110[21:0]} ;
    wire [22:0] sum128_64_wire56  = {1'd0, sum256_128_reg111[21:0]} + {1'd0, sum256_128_reg112[21:0]} ;
    wire [22:0] sum128_64_wire57  = {1'd0, sum256_128_reg113[21:0]} + {1'd0, sum256_128_reg114[21:0]} ;
    wire [22:0] sum128_64_wire58  = {1'd0, sum256_128_reg115[21:0]} + {1'd0, sum256_128_reg116[21:0]} ;
    wire [22:0] sum128_64_wire59  = {1'd0, sum256_128_reg117[21:0]} + {1'd0, sum256_128_reg118[21:0]} ;
    wire [22:0] sum128_64_wire60  = {1'd0, sum256_128_reg119[21:0]} + {1'd0, sum256_128_reg120[21:0]} ;
    wire [22:0] sum128_64_wire61  = {1'd0, sum256_128_reg121[21:0]} + {1'd0, sum256_128_reg122[21:0]} ;
    wire [22:0] sum128_64_wire62  = {1'd0, sum256_128_reg123[21:0]} + {1'd0, sum256_128_reg124[21:0]} ;
    wire [22:0] sum128_64_wire63  = {1'd0, sum256_128_reg125[21:0]} + {1'd0, sum256_128_reg126[21:0]} ;
    wire [22:0] sum128_64_wire64  = {1'd0, sum256_128_reg127[21:0]} + {1'd0, sum256_128_reg128[21:0]} ;
							
    wire [23:0] sum64_32_wire01 = {1'd0, sum128_64_wire01[22:0]} + {1'd0, sum128_64_wire02[22:0]} ;
    wire [23:0] sum64_32_wire02 = {1'd0, sum128_64_wire03[22:0]} + {1'd0, sum128_64_wire04[22:0]} ;
    wire [23:0] sum64_32_wire03 = {1'd0, sum128_64_wire05[22:0]} + {1'd0, sum128_64_wire06[22:0]} ;
    wire [23:0] sum64_32_wire04 = {1'd0, sum128_64_wire07[22:0]} + {1'd0, sum128_64_wire08[22:0]} ;
    wire [23:0] sum64_32_wire05 = {1'd0, sum128_64_wire09[22:0]} + {1'd0, sum128_64_wire10[22:0]} ;
    wire [23:0] sum64_32_wire06 = {1'd0, sum128_64_wire11[22:0]} + {1'd0, sum128_64_wire12[22:0]} ;
    wire [23:0] sum64_32_wire07 = {1'd0, sum128_64_wire13[22:0]} + {1'd0, sum128_64_wire14[22:0]} ;
    wire [23:0] sum64_32_wire08 = {1'd0, sum128_64_wire15[22:0]} + {1'd0, sum128_64_wire16[22:0]} ;
    wire [23:0] sum64_32_wire09 = {1'd0, sum128_64_wire17[22:0]} + {1'd0, sum128_64_wire18[22:0]} ;
    wire [23:0] sum64_32_wire10 = {1'd0, sum128_64_wire19[22:0]} + {1'd0, sum128_64_wire20[22:0]} ;
    wire [23:0] sum64_32_wire11 = {1'd0, sum128_64_wire21[22:0]} + {1'd0, sum128_64_wire22[22:0]} ;
    wire [23:0] sum64_32_wire12 = {1'd0, sum128_64_wire23[22:0]} + {1'd0, sum128_64_wire24[22:0]} ;
    wire [23:0] sum64_32_wire13 = {1'd0, sum128_64_wire25[22:0]} + {1'd0, sum128_64_wire26[22:0]} ;
    wire [23:0] sum64_32_wire14 = {1'd0, sum128_64_wire27[22:0]} + {1'd0, sum128_64_wire28[22:0]} ;
    wire [23:0] sum64_32_wire15 = {1'd0, sum128_64_wire29[22:0]} + {1'd0, sum128_64_wire30[22:0]} ;
    wire [23:0] sum64_32_wire16 = {1'd0, sum128_64_wire31[22:0]} + {1'd0, sum128_64_wire32[22:0]} ;
    wire [23:0] sum64_32_wire17 = {1'd0, sum128_64_wire33[22:0]} + {1'd0, sum128_64_wire34[22:0]} ;
    wire [23:0] sum64_32_wire18 = {1'd0, sum128_64_wire35[22:0]} + {1'd0, sum128_64_wire36[22:0]} ;
    wire [23:0] sum64_32_wire19 = {1'd0, sum128_64_wire37[22:0]} + {1'd0, sum128_64_wire38[22:0]} ;
    wire [23:0] sum64_32_wire20 = {1'd0, sum128_64_wire39[22:0]} + {1'd0, sum128_64_wire40[22:0]} ;
    wire [23:0] sum64_32_wire21 = {1'd0, sum128_64_wire41[22:0]} + {1'd0, sum128_64_wire42[22:0]} ;
    wire [23:0] sum64_32_wire22 = {1'd0, sum128_64_wire43[22:0]} + {1'd0, sum128_64_wire44[22:0]} ;
    wire [23:0] sum64_32_wire23 = {1'd0, sum128_64_wire45[22:0]} + {1'd0, sum128_64_wire46[22:0]} ;
    wire [23:0] sum64_32_wire24 = {1'd0, sum128_64_wire47[22:0]} + {1'd0, sum128_64_wire48[22:0]} ;
    wire [23:0] sum64_32_wire25 = {1'd0, sum128_64_wire49[22:0]} + {1'd0, sum128_64_wire50[22:0]} ;
    wire [23:0] sum64_32_wire26 = {1'd0, sum128_64_wire51[22:0]} + {1'd0, sum128_64_wire52[22:0]} ;
    wire [23:0] sum64_32_wire27 = {1'd0, sum128_64_wire53[22:0]} + {1'd0, sum128_64_wire54[22:0]} ;
    wire [23:0] sum64_32_wire28 = {1'd0, sum128_64_wire55[22:0]} + {1'd0, sum128_64_wire56[22:0]} ;
    wire [23:0] sum64_32_wire29 = {1'd0, sum128_64_wire57[22:0]} + {1'd0, sum128_64_wire58[22:0]} ;
    wire [23:0] sum64_32_wire30 = {1'd0, sum128_64_wire59[22:0]} + {1'd0, sum128_64_wire60[22:0]} ;
    wire [23:0] sum64_32_wire31 = {1'd0, sum128_64_wire61[22:0]} + {1'd0, sum128_64_wire62[22:0]} ;
    wire [23:0] sum64_32_wire32 = {1'd0, sum128_64_wire63[22:0]} + {1'd0, sum128_64_wire64[22:0]} ;

	
    reg [23:0] sum64_32_reg01, sum64_32_reg02, sum64_32_reg03, sum64_32_reg04,
                sum64_32_reg05, sum64_32_reg06, sum64_32_reg07, sum64_32_reg08,
                sum64_32_reg09, sum64_32_reg10, sum64_32_reg11, sum64_32_reg12,
                sum64_32_reg13, sum64_32_reg14, sum64_32_reg15, sum64_32_reg16,
                sum64_32_reg17, sum64_32_reg18, sum64_32_reg19, sum64_32_reg20,
                sum64_32_reg21, sum64_32_reg22, sum64_32_reg23, sum64_32_reg24,
                sum64_32_reg25, sum64_32_reg26, sum64_32_reg27, sum64_32_reg28,
                sum64_32_reg29, sum64_32_reg30, sum64_32_reg31, sum64_32_reg32;
	
    always @ (posedge clk) begin
		if(rst) begin
            sum64_32_reg01[23:0] <= #DLY 24'd0 ;
            sum64_32_reg02[23:0] <= #DLY 24'd0 ;
            sum64_32_reg03[23:0] <= #DLY 24'd0 ;
            sum64_32_reg04[23:0] <= #DLY 24'd0 ;
            sum64_32_reg05[23:0] <= #DLY 24'd0 ;
            sum64_32_reg06[23:0] <= #DLY 24'd0 ;
            sum64_32_reg07[23:0] <= #DLY 24'd0 ;
            sum64_32_reg08[23:0] <= #DLY 24'd0 ;
            sum64_32_reg09[23:0] <= #DLY 24'd0 ;
            sum64_32_reg10[23:0] <= #DLY 24'd0 ;
            sum64_32_reg11[23:0] <= #DLY 24'd0 ;
            sum64_32_reg12[23:0] <= #DLY 24'd0 ;
            sum64_32_reg13[23:0] <= #DLY 24'd0 ;
            sum64_32_reg14[23:0] <= #DLY 24'd0 ;
            sum64_32_reg15[23:0] <= #DLY 24'd0 ;
            sum64_32_reg16[23:0] <= #DLY 24'd0 ;
            sum64_32_reg17[23:0] <= #DLY 24'd0 ;
            sum64_32_reg18[23:0] <= #DLY 24'd0 ;
            sum64_32_reg19[23:0] <= #DLY 24'd0 ;
            sum64_32_reg20[23:0] <= #DLY 24'd0 ;
            sum64_32_reg21[23:0] <= #DLY 24'd0 ;
            sum64_32_reg22[23:0] <= #DLY 24'd0 ;
            sum64_32_reg23[23:0] <= #DLY 24'd0 ;
            sum64_32_reg24[23:0] <= #DLY 24'd0 ;
            sum64_32_reg25[23:0] <= #DLY 24'd0 ;
            sum64_32_reg26[23:0] <= #DLY 24'd0 ;
            sum64_32_reg27[23:0] <= #DLY 24'd0 ;
            sum64_32_reg28[23:0] <= #DLY 24'd0 ;
            sum64_32_reg29[23:0] <= #DLY 24'd0 ;
            sum64_32_reg30[23:0] <= #DLY 24'd0 ;
            sum64_32_reg31[23:0] <= #DLY 24'd0 ;
            sum64_32_reg32[23:0] <= #DLY 24'd0 ;
		end else begin
            sum64_32_reg01[23:0] <= #DLY sum64_32_wire01[23:0] ;
            sum64_32_reg02[23:0] <= #DLY sum64_32_wire02[23:0] ;
            sum64_32_reg03[23:0] <= #DLY sum64_32_wire03[23:0] ;
            sum64_32_reg04[23:0] <= #DLY sum64_32_wire04[23:0] ;
            sum64_32_reg05[23:0] <= #DLY sum64_32_wire05[23:0] ;
            sum64_32_reg06[23:0] <= #DLY sum64_32_wire06[23:0] ;
            sum64_32_reg07[23:0] <= #DLY sum64_32_wire07[23:0] ;
            sum64_32_reg08[23:0] <= #DLY sum64_32_wire08[23:0] ;
            sum64_32_reg09[23:0] <= #DLY sum64_32_wire09[23:0] ;
            sum64_32_reg10[23:0] <= #DLY sum64_32_wire10[23:0] ;
            sum64_32_reg11[23:0] <= #DLY sum64_32_wire11[23:0] ;
            sum64_32_reg12[23:0] <= #DLY sum64_32_wire12[23:0] ;
            sum64_32_reg13[23:0] <= #DLY sum64_32_wire13[23:0] ;
            sum64_32_reg14[23:0] <= #DLY sum64_32_wire14[23:0] ;
            sum64_32_reg15[23:0] <= #DLY sum64_32_wire15[23:0] ;
            sum64_32_reg16[23:0] <= #DLY sum64_32_wire16[23:0] ;
            sum64_32_reg17[23:0] <= #DLY sum64_32_wire17[23:0] ;
            sum64_32_reg18[23:0] <= #DLY sum64_32_wire18[23:0] ;
            sum64_32_reg19[23:0] <= #DLY sum64_32_wire19[23:0] ;
            sum64_32_reg20[23:0] <= #DLY sum64_32_wire20[23:0] ;
            sum64_32_reg21[23:0] <= #DLY sum64_32_wire21[23:0] ;
            sum64_32_reg22[23:0] <= #DLY sum64_32_wire22[23:0] ;
            sum64_32_reg23[23:0] <= #DLY sum64_32_wire23[23:0] ;
            sum64_32_reg24[23:0] <= #DLY sum64_32_wire24[23:0] ;
            sum64_32_reg25[23:0] <= #DLY sum64_32_wire25[23:0] ;
            sum64_32_reg26[23:0] <= #DLY sum64_32_wire26[23:0] ;
            sum64_32_reg27[23:0] <= #DLY sum64_32_wire27[23:0] ;
            sum64_32_reg28[23:0] <= #DLY sum64_32_wire28[23:0] ;
            sum64_32_reg29[23:0] <= #DLY sum64_32_wire29[23:0] ;
            sum64_32_reg30[23:0] <= #DLY sum64_32_wire30[23:0] ;
            sum64_32_reg31[23:0] <= #DLY sum64_32_wire31[23:0] ;
            sum64_32_reg32[23:0] <= #DLY sum64_32_wire32[23:0] ;
		end
	end

    /****************************
    // pipeline[36] Active
    ****************************/
    wire [24:0] sum32_16_wire01 = {1'd0, sum64_32_reg01[23:0]} + {1'd0, sum64_32_reg02[23:0]} ;
    wire [24:0] sum32_16_wire02 = {1'd0, sum64_32_reg03[23:0]} + {1'd0, sum64_32_reg04[23:0]} ;
    wire [24:0] sum32_16_wire03 = {1'd0, sum64_32_reg05[23:0]} + {1'd0, sum64_32_reg06[23:0]} ;
    wire [24:0] sum32_16_wire04 = {1'd0, sum64_32_reg07[23:0]} + {1'd0, sum64_32_reg08[23:0]} ;
    wire [24:0] sum32_16_wire05 = {1'd0, sum64_32_reg09[23:0]} + {1'd0, sum64_32_reg10[23:0]} ;
    wire [24:0] sum32_16_wire06 = {1'd0, sum64_32_reg11[23:0]} + {1'd0, sum64_32_reg12[23:0]} ;
    wire [24:0] sum32_16_wire07 = {1'd0, sum64_32_reg13[23:0]} + {1'd0, sum64_32_reg14[23:0]} ;
    wire [24:0] sum32_16_wire08 = {1'd0, sum64_32_reg15[23:0]} + {1'd0, sum64_32_reg16[23:0]} ;
    wire [24:0] sum32_16_wire09 = {1'd0, sum64_32_reg17[23:0]} + {1'd0, sum64_32_reg18[23:0]} ;
    wire [24:0] sum32_16_wire10 = {1'd0, sum64_32_reg19[23:0]} + {1'd0, sum64_32_reg20[23:0]} ;
    wire [24:0] sum32_16_wire11 = {1'd0, sum64_32_reg21[23:0]} + {1'd0, sum64_32_reg22[23:0]} ;
    wire [24:0] sum32_16_wire12 = {1'd0, sum64_32_reg23[23:0]} + {1'd0, sum64_32_reg24[23:0]} ;
    wire [24:0] sum32_16_wire13 = {1'd0, sum64_32_reg25[23:0]} + {1'd0, sum64_32_reg26[23:0]} ;
    wire [24:0] sum32_16_wire14 = {1'd0, sum64_32_reg27[23:0]} + {1'd0, sum64_32_reg28[23:0]} ;
    wire [24:0] sum32_16_wire15 = {1'd0, sum64_32_reg29[23:0]} + {1'd0, sum64_32_reg30[23:0]} ;
    wire [24:0] sum32_16_wire16 = {1'd0, sum64_32_reg31[23:0]} + {1'd0, sum64_32_reg32[23:0]} ;

    wire [25:0] sum16_8_wire01 = {1'd0, sum32_16_wire01[24:0]} + {1'd0, sum32_16_wire02[24:0]} ;
    wire [25:0] sum16_8_wire02 = {1'd0, sum32_16_wire03[24:0]} + {1'd0, sum32_16_wire04[24:0]} ;
    wire [25:0] sum16_8_wire03 = {1'd0, sum32_16_wire05[24:0]} + {1'd0, sum32_16_wire06[24:0]} ;
    wire [25:0] sum16_8_wire04 = {1'd0, sum32_16_wire07[24:0]} + {1'd0, sum32_16_wire08[24:0]} ;
    wire [25:0] sum16_8_wire05 = {1'd0, sum32_16_wire09[24:0]} + {1'd0, sum32_16_wire10[24:0]} ;
    wire [25:0] sum16_8_wire06 = {1'd0, sum32_16_wire11[24:0]} + {1'd0, sum32_16_wire12[24:0]} ;
    wire [25:0] sum16_8_wire07 = {1'd0, sum32_16_wire13[24:0]} + {1'd0, sum32_16_wire14[24:0]} ;
    wire [25:0] sum16_8_wire08 = {1'd0, sum32_16_wire15[24:0]} + {1'd0, sum32_16_wire16[24:0]} ;

	reg [25:0] sum16_8_reg01, sum16_8_reg02, sum16_8_reg03, sum16_8_reg04,
               sum16_8_reg05, sum16_8_reg06, sum16_8_reg07, sum16_8_reg08;

    always @ (posedge clk) begin
		if(rst) begin
		    sum16_8_reg01[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg02[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg03[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg04[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg05[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg06[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg07[25:0] <= #DLY 26'd0 ;
		    sum16_8_reg08[25:0] <= #DLY 26'd0 ;
		end else begin
		    sum16_8_reg01[25:0] <= #DLY sum16_8_wire01[25:0] ;
		    sum16_8_reg02[25:0] <= #DLY sum16_8_wire02[25:0] ;
		    sum16_8_reg03[25:0] <= #DLY sum16_8_wire03[25:0] ;
		    sum16_8_reg04[25:0] <= #DLY sum16_8_wire04[25:0] ;
		    sum16_8_reg05[25:0] <= #DLY sum16_8_wire05[25:0] ;
		    sum16_8_reg06[25:0] <= #DLY sum16_8_wire06[25:0] ;
		    sum16_8_reg07[25:0] <= #DLY sum16_8_wire07[25:0] ;
		    sum16_8_reg08[25:0] <= #DLY sum16_8_wire08[25:0] ;
		end
	end
  
    /****************************
    // pipeline[37] Active
    ****************************/
    wire [26:0] sum8_4_wire01 = {1'd0, sum16_8_reg01[25:0]} + {1'd0, sum16_8_reg02[25:0]} ;
    wire [26:0] sum8_4_wire02 = {1'd0, sum16_8_reg03[25:0]} + {1'd0, sum16_8_reg04[25:0]} ;
    wire [26:0] sum8_4_wire03 = {1'd0, sum16_8_reg05[25:0]} + {1'd0, sum16_8_reg06[25:0]} ;
    wire [26:0] sum8_4_wire04 = {1'd0, sum16_8_reg07[25:0]} + {1'd0, sum16_8_reg08[25:0]} ;
	
    wire [27:0] sum4_2_wire01 = {1'd0, sum8_4_wire01[26:0]} + {1'd0, sum8_4_wire02[26:0]} ;
    wire [27:0] sum4_2_wire02 = {1'd0, sum8_4_wire03[26:0]} + {1'd0, sum8_4_wire04[26:0]} ;
	
	reg [27:0] sum4_2_reg01, sum4_2_reg02 ;
	
    always @ (posedge clk) begin
		if(rst) begin
		    sum4_2_reg01[27:0] <= #DLY 28'd0 ;
		    sum4_2_reg02[27:0] <= #DLY 28'd0 ;
		end else begin
		    sum4_2_reg01[27:0] <= #DLY sum4_2_wire01[27:0] ;
		    sum4_2_reg02[27:0] <= #DLY sum4_2_wire02[27:0] ;
		end
	end
  
    /****************************
    // pipeline[38] Active
    ****************************/
    wire [28:0] sum1_wire = {1'd0, sum4_2_reg01[27:0]} + {1'd0, sum4_2_reg02[27:0]} ;
    reg  [28:0] sum1_reg;

    always @ (posedge clk) begin
		if(rst) begin
			sum1_reg[28:0] <= #DLY 29'd0 ;
		end else begin
			sum1_reg[28:0] <= #DLY sum1_wire[28:0] ;
		end
	end
	
    /****************************
    // pipeline[39] Active
    ****************************/
    reg  [29:0] sum_reg00, sum_reg01, sum_reg02, sum_reg03,
                sum_reg04, sum_reg05, sum_reg06, sum_reg07,
                sum_reg08, sum_reg09, sum_reg10, sum_reg11,
                sum_reg12, sum_reg13, sum_reg14, sum_reg15,
                sum_reg16, sum_reg17, sum_reg18, sum_reg19,
                sum_reg20, sum_reg21, sum_reg22, sum_reg23,
                sum_reg24, sum_reg25, sum_reg26, sum_reg27,
                sum_reg28, sum_reg29, sum_reg30, sum_reg31;

    always @ (posedge clk) begin
		if(rst) begin
			sum_reg00[29:0] <= #DLY 30'd0 ;
			sum_reg01[29:0] <= #DLY 30'd0 ;
			sum_reg02[29:0] <= #DLY 30'd0 ;
			sum_reg03[29:0] <= #DLY 30'd0 ;
			sum_reg04[29:0] <= #DLY 30'd0 ;
			sum_reg05[29:0] <= #DLY 30'd0 ;
			sum_reg06[29:0] <= #DLY 30'd0 ;
			sum_reg07[29:0] <= #DLY 30'd0 ;
			sum_reg08[29:0] <= #DLY 30'd0 ;
			sum_reg09[29:0] <= #DLY 30'd0 ;
			sum_reg10[29:0] <= #DLY 30'd0 ;
			sum_reg11[29:0] <= #DLY 30'd0 ;
			sum_reg12[29:0] <= #DLY 30'd0 ;
			sum_reg13[29:0] <= #DLY 30'd0 ;
			sum_reg14[29:0] <= #DLY 30'd0 ;
			sum_reg15[29:0] <= #DLY 30'd0 ;
			sum_reg16[29:0] <= #DLY 30'd0 ;
			sum_reg17[29:0] <= #DLY 30'd0 ;
			sum_reg18[29:0] <= #DLY 30'd0 ;
			sum_reg19[29:0] <= #DLY 30'd0 ;
			sum_reg20[29:0] <= #DLY 30'd0 ;
			sum_reg21[29:0] <= #DLY 30'd0 ;
			sum_reg22[29:0] <= #DLY 30'd0 ;
			sum_reg23[29:0] <= #DLY 30'd0 ;
			sum_reg24[29:0] <= #DLY 30'd0 ;
			sum_reg25[29:0] <= #DLY 30'd0 ;
			sum_reg26[29:0] <= #DLY 30'd0 ;
			sum_reg27[29:0] <= #DLY 30'd0 ;
			sum_reg28[29:0] <= #DLY 30'd0 ;
			sum_reg29[29:0] <= #DLY 30'd0 ;
			sum_reg30[29:0] <= #DLY 30'd0 ;
			sum_reg31[29:0] <= #DLY 30'd0 ;
		end else if(~loop_flg_hld[39] & loop_flg_hld[40]) begin
			sum_reg00[29:0] <= #DLY {1'd0, sum1_reg[28:0]} ;
			sum_reg01[29:0] <= #DLY 30'd0 ;
			sum_reg02[29:0] <= #DLY 30'd0 ;
			sum_reg03[29:0] <= #DLY 30'd0 ;
			sum_reg04[29:0] <= #DLY 30'd0 ;
			sum_reg05[29:0] <= #DLY 30'd0 ;
			sum_reg06[29:0] <= #DLY 30'd0 ;
			sum_reg07[29:0] <= #DLY 30'd0 ;
			sum_reg08[29:0] <= #DLY 30'd0 ;
			sum_reg09[29:0] <= #DLY 30'd0 ;
			sum_reg10[29:0] <= #DLY 30'd0 ;
			sum_reg11[29:0] <= #DLY 30'd0 ;
			sum_reg12[29:0] <= #DLY 30'd0 ;
			sum_reg13[29:0] <= #DLY 30'd0 ;
			sum_reg14[29:0] <= #DLY 30'd0 ;
			sum_reg15[29:0] <= #DLY 30'd0 ;
			sum_reg16[29:0] <= #DLY 30'd0 ;
			sum_reg17[29:0] <= #DLY 30'd0 ;
			sum_reg18[29:0] <= #DLY 30'd0 ;
			sum_reg19[29:0] <= #DLY 30'd0 ;
			sum_reg20[29:0] <= #DLY 30'd0 ;
			sum_reg21[29:0] <= #DLY 30'd0 ;
			sum_reg22[29:0] <= #DLY 30'd0 ;
			sum_reg23[29:0] <= #DLY 30'd0 ;
			sum_reg24[29:0] <= #DLY 30'd0 ;
			sum_reg25[29:0] <= #DLY 30'd0 ;
			sum_reg26[29:0] <= #DLY 30'd0 ;
			sum_reg27[29:0] <= #DLY 30'd0 ;
			sum_reg28[29:0] <= #DLY 30'd0 ;
			sum_reg29[29:0] <= #DLY 30'd0 ;
			sum_reg30[29:0] <= #DLY 30'd0 ;
			sum_reg31[29:0] <= #DLY 30'd0 ;
		end else if(pipeline_cnt[39]) begin
			if(cyc32_cnt_dd39[5:0] ==  6'd0) sum_reg00[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg00[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd1) sum_reg01[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg01[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd2) sum_reg02[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg02[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd3) sum_reg03[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg03[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd4) sum_reg04[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg04[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd5) sum_reg05[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg05[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd6) sum_reg06[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg06[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd7) sum_reg07[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg07[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd8) sum_reg08[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg08[29:0] ;
			if(cyc32_cnt_dd39[5:0] ==  6'd9) sum_reg09[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg09[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd10) sum_reg10[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg10[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd11) sum_reg11[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg11[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd12) sum_reg12[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg12[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd13) sum_reg13[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg13[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd14) sum_reg14[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg14[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd15) sum_reg15[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg15[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd16) sum_reg16[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg16[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd17) sum_reg17[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg17[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd18) sum_reg18[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg18[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd19) sum_reg19[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg19[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd20) sum_reg20[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg20[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd21) sum_reg21[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg21[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd22) sum_reg22[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg22[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd23) sum_reg23[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg23[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd24) sum_reg24[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg24[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd25) sum_reg25[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg25[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd26) sum_reg26[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg26[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd27) sum_reg27[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg27[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd28) sum_reg28[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg28[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd29) sum_reg29[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg29[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd30) sum_reg30[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg30[29:0] ;
			if(cyc32_cnt_dd39[5:0] == 6'd31) sum_reg31[29:0] <= #DLY {1'd0, sum1_reg[28:0]} + sum_reg31[29:0] ;
		end
	end


    /****************************
    // pipeline[40] Active
    ****************************/
	assign out_en  = (pipeline_cnt[40] & loop_flg_hld[40]);
	assign out_dat[19:0] = (cyc32_cnt_dd40[5:0] ==  6'd0)? sum_reg00[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd1)? sum_reg01[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd2)? sum_reg02[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd3)? sum_reg03[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd4)? sum_reg04[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd5)? sum_reg05[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd6)? sum_reg06[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd7)? sum_reg07[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd8)? sum_reg08[29:10] :
                           (cyc32_cnt_dd40[5:0] ==  6'd9)? sum_reg09[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd10)? sum_reg10[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd11)? sum_reg11[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd12)? sum_reg12[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd13)? sum_reg13[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd14)? sum_reg14[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd15)? sum_reg15[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd16)? sum_reg16[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd17)? sum_reg17[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd18)? sum_reg18[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd19)? sum_reg19[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd20)? sum_reg20[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd21)? sum_reg21[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd22)? sum_reg22[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd23)? sum_reg23[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd24)? sum_reg24[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd25)? sum_reg25[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd26)? sum_reg26[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd27)? sum_reg27[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd28)? sum_reg28[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd29)? sum_reg29[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd30)? sum_reg30[29:10] :
                           (cyc32_cnt_dd40[5:0] == 6'd31)? sum_reg31[29:10] : 20'd0 ;

endmodule
